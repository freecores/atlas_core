-- ########################################################
-- #         << ATLAS Project - Bootloader ROM >>         #
-- # **************************************************** #
-- #  2kB ROM initialized with Atlas-2k bootloader.       #
-- # **************************************************** #
-- #  Last modified: 04.05.2014                           #
-- # **************************************************** #
-- #  by Stephan Nolting 4788, Hanover, Germany           #
-- ########################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.atlas_core_package.all;

entity BOOT_MEM is
	port	(
				-- Host Interface --
				CLK_I           : in  std_logic; -- global clock line
				I_ADR_I         : in  std_logic_vector(15 downto 0); -- instruction adr
				I_EN_I          : in  std_logic; -- IR update
				I_DAT_O         : out std_logic_vector(15 downto 0); -- instruction out
				D_EN_I          : in  std_logic; -- access enable
				D_RW_I          : in  std_logic; -- read/write
				D_ADR_I         : in  std_logic_vector(15 downto 0); -- data adr
				D_DAT_I         : in  std_logic_vector(15 downto 0); -- data in
				D_DAT_O         : out std_logic_vector(15 downto 0)  -- data out
			);
end BOOT_MEM;

architecture BOOT_MEM_STRUCTURE of BOOT_MEM is

	-- Internal constants(configuration --
	constant mem_size_c      : natural := 2048; -- 2kB
	constant log2_mem_size_c : natural := log2(mem_size_c/2); -- address width (word boundary!)

	-- Memory Type --
	type mem_file_t is array (0 to (mem_size_c/2)-1) of std_logic_vector(15 downto 0); -- word mem!

	-- MEMORY IMAGE (Bootloader Program) --
	------------------------------------------------------
	constant BOOT_MEM_FILE_C : mem_file_t :=
    (
		000000 => x"bc0e", -- B
		000001 => x"bc04", -- B
		000002 => x"bc03", -- B
		000003 => x"bc02", -- B
		000004 => x"bc01", -- B
		000005 => x"c000", -- LDIL
		000006 => x"cc00", -- LDIH
		000007 => x"ec8a", -- MCR
		000008 => x"cc19", -- LDIH
		000009 => x"ed0f", -- MCR
		000010 => x"c528", -- LDIL
		000011 => x"c907", -- LDIH
		000012 => x"be73", -- BL
		000013 => x"bc00", -- B
		000014 => x"ec11", -- MRC
		000015 => x"ec88", -- MCR
		000016 => x"ec8a", -- MCR
		000017 => x"c380", -- LDIL
		000018 => x"cff8", -- LDIH
		000019 => x"1c07", -- STSR
		000020 => x"2800", -- CLR
		000021 => x"ec08", -- MCR
		000022 => x"ec0b", -- MCR
		000023 => x"ec0d", -- MCR
		000024 => x"ec00", -- MRC
		000025 => x"ed88", -- MCR
		000026 => x"ed8b", -- MCR
		000027 => x"c064", -- LDIL
		000028 => x"ed8d", -- MCR
		000029 => x"c901", -- LDIH
		000030 => x"ed2f", -- MCR
		000031 => x"ec17", -- MRC
		000032 => x"ec97", -- MRC
		000033 => x"c160", -- LDIL
		000034 => x"c909", -- LDIH
		000035 => x"c18f", -- LDIL
		000036 => x"0923", -- ADD
		000037 => x"29b3", -- CLR
		000038 => x"2a44", -- CLR
		000039 => x"100a", -- SUBS
		000040 => x"149b", -- SBCS
		000041 => x"9003", -- BMI
		000042 => x"0241", -- INC
		000043 => x"bdfc", -- B
		000044 => x"ed49", -- MCR
		000045 => x"ec22", -- MRC
		000046 => x"d406", -- SBR
		000047 => x"ed0a", -- MCR
		000048 => x"c53c", -- LDIL
		000049 => x"c905", -- LDIH
		000050 => x"be4d", -- BL
		000051 => x"c132", -- LDIL
		000052 => x"c906", -- LDIH
		000053 => x"be4a", -- BL
		000054 => x"ee11", -- MRC
		000055 => x"be4c", -- BL
		000056 => x"c142", -- LDIL
		000057 => x"c906", -- LDIH
		000058 => x"be45", -- BL
		000059 => x"ee97", -- MRC
		000060 => x"ee17", -- MRC
		000061 => x"be46", -- BL
		000062 => x"0250", -- MOV
		000063 => x"be44", -- BL
		000064 => x"be40", -- BL
		000065 => x"ec27", -- MRC
		000066 => x"c083", -- LDIL
		000067 => x"2001", -- AND
		000068 => x"c330", -- LDIL
		000069 => x"0b60", -- ADD
		000070 => x"bc0f", -- B
		000071 => x"c55a", -- LDIL
		000072 => x"c906", -- LDIH
		000073 => x"be36", -- BL
		000074 => x"c14c", -- LDIL
		000075 => x"c907", -- LDIH
		000076 => x"be33", -- BL
		000077 => x"c512", -- LDIL
		000078 => x"c907", -- LDIH
		000079 => x"be30", -- BL
		000080 => x"be32", -- BL
		000081 => x"0300", -- MOV
		000082 => x"0080", -- MOV
		000083 => x"be2e", -- BL
		000084 => x"be2c", -- BL
		000085 => x"c0b0", -- LDIL
		000086 => x"181e", -- CMP
		000087 => x"81f0", -- BEQ
		000088 => x"c0b1", -- LDIL
		000089 => x"181e", -- CMP
		000090 => x"8085", -- BEQ
		000091 => x"c0b2", -- LDIL
		000092 => x"181e", -- CMP
		000093 => x"8052", -- BEQ
		000094 => x"c0b3", -- LDIL
		000095 => x"181e", -- CMP
		000096 => x"8019", -- BEQ
		000097 => x"c0b4", -- LDIL
		000098 => x"181e", -- CMP
		000099 => x"8021", -- BEQ
		000100 => x"c29c", -- LDIL
		000101 => x"ca83", -- LDIH
		000102 => x"c0f0", -- LDIL
		000103 => x"181e", -- CMP
		000104 => x"f705", -- RBAEQ
		000105 => x"c0e4", -- LDIL
		000106 => x"181e", -- CMP
		000107 => x"80e4", -- BEQ
		000108 => x"c2d0", -- LDIL
		000109 => x"ca85", -- LDIH
		000110 => x"c0f7", -- LDIL
		000111 => x"181e", -- CMP
		000112 => x"f705", -- RBAEQ
		000113 => x"c0f2", -- LDIL
		000114 => x"181e", -- CMP
		000115 => x"85da", -- BNE
		000116 => x"2800", -- CLR
		000117 => x"c080", -- LDIL
		000118 => x"cc80", -- LDIH
		000119 => x"ec99", -- MCR
		000120 => x"3400", -- GT
		000121 => x"c152", -- LDIL
		000122 => x"c906", -- LDIH
		000123 => x"be04", -- BL
		000124 => x"2800", -- CLR
		000125 => x"2100", -- STUB
		000126 => x"bca3", -- B
		000127 => x"bc98", -- B
		000128 => x"bc98", -- B
		000129 => x"bc98", -- B
		000130 => x"bc98", -- B
		000131 => x"bc9b", -- B
		000132 => x"c530", -- LDIL
		000133 => x"c906", -- LDIH
		000134 => x"be91", -- BL
		000135 => x"be99", -- BL
		000136 => x"edca", -- MCR
		000137 => x"be97", -- BL
		000138 => x"edc9", -- MCR
		000139 => x"c03e", -- LDIL
		000140 => x"c805", -- LDIH
		000141 => x"3404", -- GTL
		000142 => x"be8a", -- BL
		000143 => x"be90", -- BL
		000144 => x"c47e", -- LDIL
		000145 => x"cc4a", -- LDIH
		000146 => x"180e", -- CMP
		000147 => x"8489", -- BNE
		000148 => x"be8b", -- BL
		000149 => x"3f64", -- SFT
		000150 => x"2066", -- STUB
		000151 => x"be88", -- BL
		000152 => x"20e6", -- STUB
		000153 => x"be86", -- BL
		000154 => x"2166", -- STUB
		000155 => x"be84", -- BL
		000156 => x"21e6", -- STUB
		000157 => x"be82", -- BL
		000158 => x"2266", -- STUB
		000159 => x"be80", -- BL
		000160 => x"22e6", -- STUB
		000161 => x"be7e", -- BL
		000162 => x"2366", -- STUB
		000163 => x"c280", -- LDIL
		000164 => x"ecda", -- MCR
		000165 => x"ec5e", -- MCR
		000166 => x"be79", -- BL
		000167 => x"7f5a", -- STR
		000168 => x"ec06", -- MRC
		000169 => x"2806", -- EOR
		000170 => x"ec0e", -- MCR
		000171 => x"2400", -- LDUB
		000172 => x"1858", -- CMP
		000173 => x"85f9", -- BNE
		000174 => x"bc56", -- B
		000175 => x"c100", -- LDIL
		000176 => x"be28", -- BL
		000177 => x"c47e", -- LDIL
		000178 => x"cc4a", -- LDIH
		000179 => x"180d", -- CMP
		000180 => x"8468", -- BNE
		000181 => x"c102", -- LDIL
		000182 => x"be22", -- BL
		000183 => x"2055", -- STUB
		000184 => x"c104", -- LDIL
		000185 => x"be1f", -- BL
		000186 => x"20d5", -- STUB
		000187 => x"c106", -- LDIL
		000188 => x"be1c", -- BL
		000189 => x"2155", -- STUB
		000190 => x"c108", -- LDIL
		000191 => x"be19", -- BL
		000192 => x"21d5", -- STUB
		000193 => x"c10a", -- LDIL
		000194 => x"be16", -- BL
		000195 => x"2255", -- STUB
		000196 => x"c10c", -- LDIL
		000197 => x"be13", -- BL
		000198 => x"22d5", -- STUB
		000199 => x"c10e", -- LDIL
		000200 => x"be10", -- BL
		000201 => x"2355", -- STUB
		000202 => x"c200", -- LDIL
		000203 => x"ecca", -- MCR
		000204 => x"ec4e", -- MCR
		000205 => x"c010", -- LDIL
		000206 => x"0940", -- ADD
		000207 => x"be09", -- BL
		000208 => x"7eca", -- STR
		000209 => x"ec06", -- MRC
		000210 => x"2805", -- EOR
		000211 => x"ec0e", -- MCR
		000212 => x"2400", -- LDUB
		000213 => x"1848", -- CMP
		000214 => x"85f7", -- BNE
		000215 => x"bc2d", -- B
		000216 => x"0370", -- MOV
		000217 => x"be42", -- BL
		000218 => x"3eb0", -- SFT
		000219 => x"0121", -- INC
		000220 => x"be3f", -- BL
		000221 => x"26d3", -- ORR
		000222 => x"3460", -- RET
		000223 => x"c16a", -- LDIL
		000224 => x"c906", -- LDIH
		000225 => x"be36", -- BL
		000226 => x"be38", -- BL
		000227 => x"3c80", -- SFT
		000228 => x"be36", -- BL
		000229 => x"2490", -- ORR
		000230 => x"c47e", -- LDIL
		000231 => x"cc4a", -- LDIH
		000232 => x"1818", -- CMP
		000233 => x"8433", -- BNE
		000234 => x"be27", -- BL
		000235 => x"3c94", -- SFT
		000236 => x"2011", -- STUB
		000237 => x"be24", -- BL
		000238 => x"2091", -- STUB
		000239 => x"be22", -- BL
		000240 => x"2111", -- STUB
		000241 => x"be20", -- BL
		000242 => x"2191", -- STUB
		000243 => x"be1e", -- BL
		000244 => x"2211", -- STUB
		000245 => x"be1c", -- BL
		000246 => x"2291", -- STUB
		000247 => x"be1a", -- BL
		000248 => x"2311", -- STUB
		000249 => x"2ad5", -- CLR
		000250 => x"ecda", -- MCR
		000251 => x"ec5e", -- MCR
		000252 => x"be15", -- BL
		000253 => x"7cda", -- STR
		000254 => x"ec06", -- MRC
		000255 => x"2801", -- EOR
		000256 => x"ec0e", -- MCR
		000257 => x"2400", -- LDUB
		000258 => x"1858", -- CMP
		000259 => x"85f9", -- BNE
		000260 => x"ec11", -- MRC
		000261 => x"ec8a", -- MCR
		000262 => x"c50e", -- LDIL
		000263 => x"c906", -- LDIH
		000264 => x"be0f", -- BL
		000265 => x"ec06", -- MRC
		000266 => x"2491", -- LDUB
		000267 => x"1809", -- CMP
		000268 => x"8015", -- BEQ
		000269 => x"c536", -- LDIL
		000270 => x"c907", -- LDIH
		000271 => x"be08", -- BL
		000272 => x"bccf", -- B
		000273 => x"0370", -- MOV
		000274 => x"be08", -- BL
		000275 => x"3c80", -- SFT
		000276 => x"be06", -- BL
		000277 => x"2490", -- ORR
		000278 => x"3460", -- RET
		000279 => x"bccb", -- B
		000280 => x"bcd4", -- B
		000281 => x"bcd8", -- B
		000282 => x"bcdc", -- B
		000283 => x"bc71", -- B
		000284 => x"bcc0", -- B
		000285 => x"bd30", -- B
		000286 => x"bc6f", -- B
		000287 => x"bcc2", -- B
		000288 => x"bcdb", -- B
		000289 => x"c17e", -- LDIL
		000290 => x"c906", -- LDIH
		000291 => x"bebf", -- BL
		000292 => x"24aa", -- LDUBS
		000293 => x"8016", -- BEQ
		000294 => x"c0a2", -- LDIL
		000295 => x"beca", -- BL
		000296 => x"24a2", -- LDUB
		000297 => x"be20", -- BL
		000298 => x"24b3", -- LDUB
		000299 => x"be1e", -- BL
		000300 => x"24c4", -- LDUB
		000301 => x"be1c", -- BL
		000302 => x"24d5", -- LDUB
		000303 => x"be1a", -- BL
		000304 => x"24e6", -- LDUB
		000305 => x"be18", -- BL
		000306 => x"c0a2", -- LDIL
		000307 => x"bebe", -- BL
		000308 => x"beb8", -- BL
		000309 => x"c54e", -- LDIL
		000310 => x"c906", -- LDIH
		000311 => x"beab", -- BL
		000312 => x"ee06", -- MRC
		000313 => x"bee7", -- BL
		000314 => x"beb2", -- BL
		000315 => x"beb1", -- BL
		000316 => x"beb0", -- BL
		000317 => x"beaf", -- BL
		000318 => x"c080", -- LDIL
		000319 => x"ccc0", -- LDIH
		000320 => x"1c01", -- STSR
		000321 => x"2800", -- CLR
		000322 => x"ed0f", -- MCR
		000323 => x"ec88", -- MCR
		000324 => x"ec8b", -- MCR
		000325 => x"ec8c", -- MCR
		000326 => x"ec8a", -- MCR
		000327 => x"ec89", -- MCR
		000328 => x"3400", -- GT
		000329 => x"0370", -- MOV
		000330 => x"3c90", -- SFT
		000331 => x"bea6", -- BL
		000332 => x"3c90", -- SFT
		000333 => x"bea4", -- BL
		000334 => x"3460", -- RET
		000335 => x"c522", -- LDIL
		000336 => x"c906", -- LDIH
		000337 => x"be91", -- BL
		000338 => x"bea9", -- BL
		000339 => x"c13e", -- LDIL
		000340 => x"c905", -- LDIH
		000341 => x"3424", -- GTL
		000342 => x"ecca", -- MCR
		000343 => x"be95", -- BL
		000344 => x"c280", -- LDIL
		000345 => x"c00f", -- LDIL
		000346 => x"2058", -- ANDS
		000347 => x"840e", -- BNE
		000348 => x"be90", -- BL
		000349 => x"c0a4", -- LDIL
		000350 => x"be93", -- BL
		000351 => x"ee12", -- MRC
		000352 => x"bec0", -- BL
		000353 => x"c0ae", -- LDIL
		000354 => x"be8f", -- BL
		000355 => x"0250", -- MOV
		000356 => x"bebc", -- BL
		000357 => x"c0ba", -- LDIL
		000358 => x"be8b", -- BL
		000359 => x"c0a0", -- LDIL
		000360 => x"be89", -- BL
		000361 => x"7a5a", -- LDR
		000362 => x"c0a0", -- LDIL
		000363 => x"be86", -- BL
		000364 => x"beb4", -- BL
		000365 => x"c00f", -- LDIL
		000366 => x"2058", -- ANDS
		000367 => x"8414", -- BNE
		000368 => x"c0a0", -- LDIL
		000369 => x"be80", -- BL
		000370 => x"be7f", -- BL
		000371 => x"c010", -- LDIL
		000372 => x"1250", -- SUB
		000373 => x"c470", -- LDIL
		000374 => x"2240", -- AND
		000375 => x"c12e", -- LDIL
		000376 => x"78c9", -- LDR
		000377 => x"3c90", -- SFT
		000378 => x"c880", -- LDIH
		000379 => x"c020", -- LDIL
		000380 => x"1818", -- CMP
		000381 => x"f8c2", -- MVHI
		000382 => x"be73", -- BL
		000383 => x"c08f", -- LDIL
		000384 => x"2014", -- AND
		000385 => x"3409", -- TEQ
		000386 => x"85f6", -- BNE
		000387 => x"ec20", -- MRC
		000388 => x"dc0f", -- STB
		000389 => x"b804", -- BTS
		000390 => x"c5fe", -- LDIL
		000391 => x"343d", -- TEQ
		000392 => x"85d1", -- BNE
		000393 => x"be6d", -- BL
		000394 => x"2800", -- CLR
		000395 => x"3400", -- GT
		000396 => x"bc54", -- B
		000397 => x"bc93", -- B
		000398 => x"c001", -- LDIL
		000399 => x"ed0c", -- MCR
		000400 => x"c050", -- LDIL
		000401 => x"c83f", -- LDIH
		000402 => x"ed0a", -- MCR
		000403 => x"c000", -- LDIL
		000404 => x"c801", -- LDIH
		000405 => x"bea9", -- BL
		000406 => x"c15c", -- LDIL
		000407 => x"c906", -- LDIH
		000408 => x"be4a", -- BL
		000409 => x"c16a", -- LDIL
		000410 => x"c906", -- LDIH
		000411 => x"be47", -- BL
		000412 => x"be5a", -- BL
		000413 => x"3c80", -- SFT
		000414 => x"be58", -- BL
		000415 => x"2410", -- ORR
		000416 => x"c4fe", -- LDIL
		000417 => x"ccca", -- LDIH
		000418 => x"1809", -- CMP
		000419 => x"8439", -- BNE
		000420 => x"c100", -- LDIL
		000421 => x"0290", -- MOV
		000422 => x"be2f", -- BL
		000423 => x"be4f", -- BL
		000424 => x"3c80", -- SFT
		000425 => x"be4d", -- BL
		000426 => x"2690", -- ORR
		000427 => x"3ed4", -- SFT
		000428 => x"2055", -- STUB
		000429 => x"c102", -- LDIL
		000430 => x"be27", -- BL
		000431 => x"be47", -- BL
		000432 => x"3c80", -- SFT
		000433 => x"be45", -- BL
		000434 => x"2690", -- ORR
		000435 => x"20d5", -- STUB
		000436 => x"c104", -- LDIL
		000437 => x"be20", -- BL
		000438 => x"c106", -- LDIL
		000439 => x"be3f", -- BL
		000440 => x"0180", -- MOV
		000441 => x"be8b", -- BL
		000442 => x"0121", -- INC
		000443 => x"c010", -- LDIL
		000444 => x"1828", -- CMP
		000445 => x"85fa", -- BNE
		000446 => x"2ad5", -- CLR
		000447 => x"be37", -- BL
		000448 => x"0180", -- MOV
		000449 => x"be83", -- BL
		000450 => x"0121", -- INC
		000451 => x"2400", -- LDUB
		000452 => x"02d1", -- INC
		000453 => x"1858", -- CMP
		000454 => x"85f9", -- BNE
		000455 => x"c001", -- LDIL
		000456 => x"ed0c", -- MCR
		000457 => x"c050", -- LDIL
		000458 => x"c83f", -- LDIH
		000459 => x"ed0a", -- MCR
		000460 => x"c00c", -- LDIL
		000461 => x"c801", -- LDIH
		000462 => x"be70", -- BL
		000463 => x"c50e", -- LDIL
		000464 => x"c906", -- LDIH
		000465 => x"be11", -- BL
		000466 => x"c68e", -- LDIL
		000467 => x"ca80", -- LDIH
		000468 => x"3450", -- GT
		000469 => x"0370", -- MOV
		000470 => x"3dd0", -- SFT
		000471 => x"be6d", -- BL
		000472 => x"0121", -- INC
		000473 => x"01d0", -- MOV
		000474 => x"be6a", -- BL
		000475 => x"3460", -- RET
		000476 => x"c51a", -- LDIL
		000477 => x"c907", -- LDIH
		000478 => x"be04", -- BL
		000479 => x"bcba", -- B
		000480 => x"bc94", -- B
		000481 => x"bca5", -- B
		000482 => x"01f0", -- MOV
		000483 => x"7829", -- LDR
		000484 => x"c080", -- LDIL
		000485 => x"ccff", -- LDIH
		000486 => x"2081", -- AND
		000487 => x"3c98", -- SFTS
		000488 => x"8003", -- BEQ
		000489 => x"be08", -- BL
		000490 => x"bdf9", -- B
		000491 => x"3430", -- RET
		000492 => x"0170", -- MOV
		000493 => x"c08d", -- LDIL
		000494 => x"be03", -- BL
		000495 => x"c08a", -- LDIL
		000496 => x"03a0", -- MOV
		000497 => x"ec22", -- MRC
		000498 => x"dc05", -- STB
		000499 => x"b9fe", -- BTS
		000500 => x"ed18", -- MCR
		000501 => x"3470", -- RET
		000502 => x"ec20", -- MRC
		000503 => x"dc8f", -- STBI
		000504 => x"b9fe", -- BTS
		000505 => x"c800", -- LDIH
		000506 => x"3470", -- RET
		000507 => x"0170", -- MOV
		000508 => x"c200", -- LDIL
		000509 => x"c184", -- LDIL
		000510 => x"bff8", -- BL
		000511 => x"c0c6", -- LDIL
		000512 => x"1809", -- CMP
		000513 => x"9003", -- BMI
		000514 => x"c0a0", -- LDIL
		000515 => x"1001", -- SUB
		000516 => x"c0b0", -- LDIL
		000517 => x"1809", -- CMP
		000518 => x"91f8", -- BMI
		000519 => x"c0c6", -- LDIL
		000520 => x"1818", -- CMP
		000521 => x"91f5", -- BMI
		000522 => x"c0b9", -- LDIL
		000523 => x"1818", -- CMP
		000524 => x"a404", -- BLS
		000525 => x"c0c1", -- LDIL
		000526 => x"1809", -- CMP
		000527 => x"a1ef", -- BHI
		000528 => x"0080", -- MOV
		000529 => x"bfe0", -- BL
		000530 => x"c030", -- LDIL
		000531 => x"1090", -- SUB
		000532 => x"c009", -- LDIL
		000533 => x"1809", -- CMP
		000534 => x"a402", -- BLS
		000535 => x"0497", -- DEC
		000536 => x"3e42", -- SFT
		000537 => x"3e42", -- SFT
		000538 => x"3e42", -- SFT
		000539 => x"3e42", -- SFT
		000540 => x"2641", -- ORR
		000541 => x"05b9", -- DECS
		000542 => x"85e0", -- BNE
		000543 => x"3420", -- RET
		000544 => x"0370", -- MOV
		000545 => x"3d42", -- SFT
		000546 => x"3d22", -- SFT
		000547 => x"3d22", -- SFT
		000548 => x"3d22", -- SFT
		000549 => x"be0f", -- BL
		000550 => x"bfcb", -- BL
		000551 => x"3d40", -- SFT
		000552 => x"be0c", -- BL
		000553 => x"bfc8", -- BL
		000554 => x"3d45", -- SFT
		000555 => x"3d25", -- SFT
		000556 => x"3d25", -- SFT
		000557 => x"3d25", -- SFT
		000558 => x"be06", -- BL
		000559 => x"bfc2", -- BL
		000560 => x"0140", -- MOV
		000561 => x"be03", -- BL
		000562 => x"bfbf", -- BL
		000563 => x"3460", -- RET
		000564 => x"c08f", -- LDIL
		000565 => x"2121", -- AND
		000566 => x"c089", -- LDIL
		000567 => x"181a", -- CMP
		000568 => x"8803", -- BCS
		000569 => x"c0b0", -- LDIL
		000570 => x"bc02", -- B
		000571 => x"c0b7", -- LDIL
		000572 => x"0892", -- ADD
		000573 => x"3470", -- RET
		000574 => x"ed0b", -- MCR
		000575 => x"ec22", -- MRC
		000576 => x"dc03", -- STB
		000577 => x"b9fe", -- BTS
		000578 => x"ec23", -- MRC
		000579 => x"3470", -- RET
		000580 => x"00f0", -- MOV
		000581 => x"c050", -- LDIL
		000582 => x"c837", -- LDIH
		000583 => x"ed0a", -- MCR
		000584 => x"c001", -- LDIL
		000585 => x"ed0c", -- MCR
		000586 => x"c006", -- LDIL
		000587 => x"bff3", -- BL
		000588 => x"c050", -- LDIL
		000589 => x"c83f", -- LDIH
		000590 => x"ed0a", -- MCR
		000591 => x"c000", -- LDIL
		000592 => x"c805", -- LDIH
		000593 => x"bfed", -- BL
		000594 => x"dc01", -- STB
		000595 => x"b805", -- BTS
		000596 => x"c546", -- LDIL
		000597 => x"c907", -- LDIH
		000598 => x"bf8c", -- BL
		000599 => x"bc42", -- B
		000600 => x"c040", -- LDIL
		000601 => x"c83f", -- LDIH
		000602 => x"ed0a", -- MCR
		000603 => x"c001", -- LDIL
		000604 => x"ed0c", -- MCR
		000605 => x"3c20", -- SFT
		000606 => x"c802", -- LDIH
		000607 => x"bfdf", -- BL
		000608 => x"03a0", -- MOV
		000609 => x"cb80", -- LDIH
		000610 => x"3ff0", -- SFT
		000611 => x"0030", -- MOV
		000612 => x"c800", -- LDIH
		000613 => x"2407", -- ORR
		000614 => x"bfd8", -- BL
		000615 => x"2800", -- CLR
		000616 => x"ed0c", -- MCR
		000617 => x"c050", -- LDIL
		000618 => x"c83f", -- LDIH
		000619 => x"ed0a", -- MCR
		000620 => x"c001", -- LDIL
		000621 => x"ed0c", -- MCR
		000622 => x"c000", -- LDIL
		000623 => x"c805", -- LDIH
		000624 => x"bfce", -- BL
		000625 => x"dc00", -- STB
		000626 => x"b9fc", -- BTS
		000627 => x"3410", -- RET
		000628 => x"00f0", -- MOV
		000629 => x"c040", -- LDIL
		000630 => x"c83f", -- LDIH
		000631 => x"ed0a", -- MCR
		000632 => x"c001", -- LDIL
		000633 => x"ed0c", -- MCR
		000634 => x"3c20", -- SFT
		000635 => x"c803", -- LDIH
		000636 => x"bfc2", -- BL
		000637 => x"0020", -- MOV
		000638 => x"c800", -- LDIH
		000639 => x"3c00", -- SFT
		000640 => x"bfbe", -- BL
		000641 => x"29b3", -- CLR
		000642 => x"ed3c", -- MCR
		000643 => x"0180", -- MOV
		000644 => x"c980", -- LDIH
		000645 => x"3410", -- RET
		000646 => x"e5b0", -- CDP
		000647 => x"ec30", -- MRC
		000648 => x"dc06", -- STB
		000649 => x"b9fe", -- BTS
		000650 => x"c306", -- LDIL
		000651 => x"200e", -- ANDS
		000652 => x"840a", -- BNE
		000653 => x"ecb1", -- MRC
		000654 => x"ef32", -- MRC
		000655 => x"2800", -- CLR
		000656 => x"009a", -- INCS
		000657 => x"0f60", -- ADC
		000658 => x"ed99", -- MCR
		000659 => x"edea", -- MCR
		000660 => x"ef34", -- MRC
		000661 => x"3470", -- RET
		000662 => x"c558", -- LDIL
		000663 => x"c907", -- LDIH
		000664 => x"bf4a", -- BL
		000665 => x"c566", -- LDIL
		000666 => x"c907", -- LDIH
		000667 => x"bf47", -- BL
		000668 => x"bf5a", -- BL
		000669 => x"2800", -- CLR
		000670 => x"3400", -- GT
		000671 => x"0170", -- MOV
		000672 => x"bf56", -- BL
		000673 => x"c08d", -- LDIL
		000674 => x"1809", -- CMP
		000675 => x"f702", -- RBAEQ
		000676 => x"c088", -- LDIL
		000677 => x"1809", -- CMP
		000678 => x"8034", -- BEQ
		000679 => x"bdf9", -- B
		000680 => x"c530", -- LDIL
		000681 => x"c906", -- LDIH
		000682 => x"bf38", -- BL
		000683 => x"bf50", -- BL
		000684 => x"edca", -- MCR
		000685 => x"bf4e", -- BL
		000686 => x"edc9", -- MCR
		000687 => x"bff0", -- BL
		000688 => x"bf3c", -- BL
		000689 => x"c53e", -- LDIL
		000690 => x"c906", -- LDIH
		000691 => x"bf2f", -- BL
		000692 => x"bf47", -- BL
		000693 => x"02c0", -- MOV
		000694 => x"bfe9", -- BL
		000695 => x"bf35", -- BL
		000696 => x"345d", -- TEQ
		000697 => x"8021", -- BEQ
		000698 => x"06d1", -- DEC
		000699 => x"bf31", -- BL
		000700 => x"c0a4", -- LDIL
		000701 => x"bf34", -- BL
		000702 => x"ee32", -- MRC
		000703 => x"bf61", -- BL
		000704 => x"ee31", -- MRC
		000705 => x"bf5f", -- BL
		000706 => x"c0ba", -- LDIL
		000707 => x"bf2e", -- BL
		000708 => x"c0a0", -- LDIL
		000709 => x"bf2c", -- BL
		000710 => x"bfc0", -- BL
		000711 => x"0260", -- MOV
		000712 => x"bf58", -- BL
		000713 => x"c320", -- LDIL
		000714 => x"c1ae", -- LDIL
		000715 => x"00e0", -- MOV
		000716 => x"bf25", -- BL
		000717 => x"3cc0", -- SFT
		000718 => x"c880", -- LDIH
		000719 => x"181e", -- CMP
		000720 => x"f8c3", -- MVHI
		000721 => x"bf20", -- BL
		000722 => x"00c0", -- MOV
		000723 => x"c880", -- LDIH
		000724 => x"181e", -- CMP
		000725 => x"f8c3", -- MVHI
		000726 => x"bf1b", -- BL
		000727 => x"eca0", -- MRC
		000728 => x"dc9f", -- STBI
		000729 => x"b9df", -- BTS
		000730 => x"bf12", -- BL
		000731 => x"c69a", -- LDIL
		000732 => x"ca80", -- LDIH
		000733 => x"3450", -- GT
		000734 => x"0d0a", -- .DW
		000735 => x"0d0a", -- .DW
		000736 => x"4174", -- .DW
		000737 => x"6c61", -- .DW
		000738 => x"732d", -- .DW
		000739 => x"324b", -- .DW
		000740 => x"2042", -- .DW
		000741 => x"6f6f", -- .DW
		000742 => x"746c", -- .DW
		000743 => x"6f61", -- .DW
		000744 => x"6465", -- .DW
		000745 => x"7220", -- .DW
		000746 => x"2d20", -- .DW
		000747 => x"5632", -- .DW
		000748 => x"3031", -- .DW
		000749 => x"3430", -- .DW
		000750 => x"3530", -- .DW
		000751 => x"340d", -- .DW
		000752 => x"0a62", -- .DW
		000753 => x"7920", -- .DW
		000754 => x"5374", -- .DW
		000755 => x"6570", -- .DW
		000756 => x"6861", -- .DW
		000757 => x"6e20", -- .DW
		000758 => x"4e6f", -- .DW
		000759 => x"6c74", -- .DW
		000760 => x"696e", -- .DW
		000761 => x"672c", -- .DW
		000762 => x"2073", -- .DW
		000763 => x"746e", -- .DW
		000764 => x"6f6c", -- .DW
		000765 => x"7469", -- .DW
		000766 => x"6e67", -- .DW
		000767 => x"4067", -- .DW
		000768 => x"6d61", -- .DW
		000769 => x"696c", -- .DW
		000770 => x"2e63", -- .DW
		000771 => x"6f6d", -- .DW
		000772 => x"0d0a", -- .DW
		000773 => x"7777", -- .DW
		000774 => x"772e", -- .DW
		000775 => x"6f70", -- .DW
		000776 => x"656e", -- .DW
		000777 => x"636f", -- .DW
		000778 => x"7265", -- .DW
		000779 => x"732e", -- .DW
		000780 => x"6f72", -- .DW
		000781 => x"672f", -- .DW
		000782 => x"7072", -- .DW
		000783 => x"6f6a", -- .DW
		000784 => x"6563", -- .DW
		000785 => x"742c", -- .DW
		000786 => x"6174", -- .DW
		000787 => x"6c61", -- .DW
		000788 => x"735f", -- .DW
		000789 => x"636f", -- .DW
		000790 => x"7265", -- .DW
		000791 => x"0d0a", -- .DW
		000792 => x"0000", -- .DW
		000793 => x"0d0a", -- .DW
		000794 => x"426f", -- .DW
		000795 => x"6f74", -- .DW
		000796 => x"2070", -- .DW
		000797 => x"6167", -- .DW
		000798 => x"653a", -- .DW
		000799 => x"2030", -- .DW
		000800 => x"7800", -- .DW
		000801 => x"0d0a", -- .DW
		000802 => x"436c", -- .DW
		000803 => x"6f63", -- .DW
		000804 => x"6b28", -- .DW
		000805 => x"487a", -- .DW
		000806 => x"293a", -- .DW
		000807 => x"2030", -- .DW
		000808 => x"7800", -- .DW
		000809 => x"426f", -- .DW
		000810 => x"6f74", -- .DW
		000811 => x"696e", -- .DW
		000812 => x"670d", -- .DW
		000813 => x"0a00", -- .DW
		000814 => x"4275", -- .DW
		000815 => x"726e", -- .DW
		000816 => x"2045", -- .DW
		000817 => x"4550", -- .DW
		000818 => x"524f", -- .DW
		000819 => x"4d0d", -- .DW
		000820 => x"0a00", -- .DW
		000821 => x"4177", -- .DW
		000822 => x"6169", -- .DW
		000823 => x"7469", -- .DW
		000824 => x"6e67", -- .DW
		000825 => x"2064", -- .DW
		000826 => x"6174", -- .DW
		000827 => x"612e", -- .DW
		000828 => x"2e2e", -- .DW
		000829 => x"0d0a", -- .DW
		000830 => x"0000", -- .DW
		000831 => x"5374", -- .DW
		000832 => x"6172", -- .DW
		000833 => x"7469", -- .DW
		000834 => x"6e67", -- .DW
		000835 => x"2069", -- .DW
		000836 => x"6d61", -- .DW
		000837 => x"6765", -- .DW
		000838 => x"2000", -- .DW
		000839 => x"446f", -- .DW
		000840 => x"776e", -- .DW
		000841 => x"6c6f", -- .DW
		000842 => x"6164", -- .DW
		000843 => x"2063", -- .DW
		000844 => x"6f6d", -- .DW
		000845 => x"706c", -- .DW
		000846 => x"6574", -- .DW
		000847 => x"650d", -- .DW
		000848 => x"0a00", -- .DW
		000849 => x"5061", -- .DW
		000850 => x"6765", -- .DW
		000851 => x"2028", -- .DW
		000852 => x"3468", -- .DW
		000853 => x"293a", -- .DW
		000854 => x"2024", -- .DW
		000855 => x"0000", -- .DW
		000856 => x"4164", -- .DW
		000857 => x"6472", -- .DW
		000858 => x"2028", -- .DW
		000859 => x"3868", -- .DW
		000860 => x"293a", -- .DW
		000861 => x"2024", -- .DW
		000862 => x"0000", -- .DW
		000863 => x"2377", -- .DW
		000864 => x"6f72", -- .DW
		000865 => x"6473", -- .DW
		000866 => x"2028", -- .DW
		000867 => x"3468", -- .DW
		000868 => x"293a", -- .DW
		000869 => x"2024", -- .DW
		000870 => x"0000", -- .DW
		000871 => x"4368", -- .DW
		000872 => x"6563", -- .DW
		000873 => x"6b73", -- .DW
		000874 => x"756d", -- .DW
		000875 => x"3a20", -- .DW
		000876 => x"2400", -- .DW
		000877 => x"0d0a", -- .DW
		000878 => x"636d", -- .DW
		000879 => x"642f", -- .DW
		000880 => x"626f", -- .DW
		000881 => x"6f74", -- .DW
		000882 => x"2d73", -- .DW
		000883 => x"7769", -- .DW
		000884 => x"7463", -- .DW
		000885 => x"683a", -- .DW
		000886 => x"0d0a", -- .DW
		000887 => x"2030", -- .DW
		000888 => x"2f27", -- .DW
		000889 => x"3030", -- .DW
		000890 => x"273a", -- .DW
		000891 => x"2028", -- .DW
		000892 => x"5265", -- .DW
		000893 => x"2d29", -- .DW
		000894 => x"5374", -- .DW
		000895 => x"6172", -- .DW
		000896 => x"7420", -- .DW
		000897 => x"636f", -- .DW
		000898 => x"6e73", -- .DW
		000899 => x"6f6c", -- .DW
		000900 => x"650d", -- .DW
		000901 => x"0a20", -- .DW
		000902 => x"312f", -- .DW
		000903 => x"2730", -- .DW
		000904 => x"3127", -- .DW
		000905 => x"3a20", -- .DW
		000906 => x"426f", -- .DW
		000907 => x"6f74", -- .DW
		000908 => x"2055", -- .DW
		000909 => x"4152", -- .DW
		000910 => x"540d", -- .DW
		000911 => x"0a20", -- .DW
		000912 => x"322f", -- .DW
		000913 => x"2731", -- .DW
		000914 => x"3027", -- .DW
		000915 => x"3a20", -- .DW
		000916 => x"426f", -- .DW
		000917 => x"6f74", -- .DW
		000918 => x"2045", -- .DW
		000919 => x"4550", -- .DW
		000920 => x"524f", -- .DW
		000921 => x"4d0d", -- .DW
		000922 => x"0a20", -- .DW
		000923 => x"332f", -- .DW
		000924 => x"2731", -- .DW
		000925 => x"3127", -- .DW
		000926 => x"3a20", -- .DW
		000927 => x"426f", -- .DW
		000928 => x"6f74", -- .DW
		000929 => x"206d", -- .DW
		000930 => x"656d", -- .DW
		000931 => x"6f72", -- .DW
		000932 => x"790d", -- .DW
		000933 => x"0a00", -- .DW
		000934 => x"2034", -- .DW
		000935 => x"3a20", -- .DW
		000936 => x"426f", -- .DW
		000937 => x"6f74", -- .DW
		000938 => x"2057", -- .DW
		000939 => x"420d", -- .DW
		000940 => x"0a20", -- .DW
		000941 => x"703a", -- .DW
		000942 => x"2042", -- .DW
		000943 => x"7572", -- .DW
		000944 => x"6e20", -- .DW
		000945 => x"4545", -- .DW
		000946 => x"5052", -- .DW
		000947 => x"4f4d", -- .DW
		000948 => x"0d0a", -- .DW
		000949 => x"2064", -- .DW
		000950 => x"3a20", -- .DW
		000951 => x"5241", -- .DW
		000952 => x"4d20", -- .DW
		000953 => x"6475", -- .DW
		000954 => x"6d70", -- .DW
		000955 => x"0d0a", -- .DW
		000956 => x"2072", -- .DW
		000957 => x"3a20", -- .DW
		000958 => x"5265", -- .DW
		000959 => x"7365", -- .DW
		000960 => x"740d", -- .DW
		000961 => x"0a20", -- .DW
		000962 => x"773a", -- .DW
		000963 => x"2057", -- .DW
		000964 => x"4220", -- .DW
		000965 => x"6475", -- .DW
		000966 => x"6d70", -- .DW
		000967 => x"0d0a", -- .DW
		000968 => x"0000", -- .DW
		000969 => x"636d", -- .DW
		000970 => x"643a", -- .DW
		000971 => x"3e20", -- .DW
		000972 => x"0000", -- .DW
		000973 => x"494d", -- .DW
		000974 => x"4147", -- .DW
		000975 => x"4520", -- .DW
		000976 => x"4552", -- .DW
		000977 => x"5221", -- .DW
		000978 => x"0d0a", -- .DW
		000979 => x"0000", -- .DW
		000980 => x"0d0a", -- .DW
		000981 => x"4952", -- .DW
		000982 => x"5120", -- .DW
		000983 => x"4552", -- .DW
		000984 => x"5221", -- .DW
		000985 => x"0d0a", -- .DW
		000986 => x"0000", -- .DW
		000987 => x"4348", -- .DW
		000988 => x"4543", -- .DW
		000989 => x"4b53", -- .DW
		000990 => x"554d", -- .DW
		000991 => x"2045", -- .DW
		000992 => x"5252", -- .DW
		000993 => x"210d", -- .DW
		000994 => x"0a00", -- .DW
		000995 => x"5350", -- .DW
		000996 => x"492f", -- .DW
		000997 => x"4545", -- .DW
		000998 => x"5052", -- .DW
		000999 => x"4f4d", -- .DW
		001000 => x"2045", -- .DW
		001001 => x"5252", -- .DW
		001002 => x"210d", -- .DW
		001003 => x"0a00", -- .DW
		001004 => x"5742", -- .DW
		001005 => x"2042", -- .DW
		001006 => x"5553", -- .DW
		001007 => x"2045", -- .DW
		001008 => x"5252", -- .DW
		001009 => x"210d", -- .DW
		001010 => x"0a00", -- .DW
		001011 => x"5072", -- .DW
		001012 => x"6573", -- .DW
		001013 => x"7320", -- .DW
		001014 => x"616e", -- .DW
		001015 => x"7920", -- .DW
		001016 => x"6b65", -- .DW
		001017 => x"790d", -- .DW
		001018 => x"0a00", -- .DW
		others => x"0000"  -- NOP
 	);
	------------------------------------------------------

begin

	-- Memory Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		MEM_FILE_ACCESS: process(CLK_I)
		begin
			if rising_edge(CLK_I) then
				-- Data Read --
				if (D_EN_I = '1') then -- valid access
					if (word_mode_en_c = true) then -- read data access
						D_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(D_ADR_I(log2_mem_size_c-1 downto 0))));
					else
						D_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(D_ADR_I(log2_mem_size_c downto 1))));
					end if;
				end if;
				-- Instruction Read --
				if (I_EN_I = '1') then
					if (word_mode_en_c = true) then
						I_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(I_ADR_I(log2_mem_size_c-1 downto 0))));
					else
						I_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(I_ADR_I(log2_mem_size_c downto 1))));
					end if;
				end if;
			end if;
		end process MEM_FILE_ACCESS;



end BOOT_MEM_STRUCTURE;
