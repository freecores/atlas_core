-- ########################################################
-- #         << ATLAS Project - Bootloader ROM >>         #
-- # **************************************************** #
-- #  Initialized with boot loader.                       #
-- # **************************************************** #
-- #  Last modified: 14.04.2014                           #
-- # **************************************************** #
-- #  by Stephan Nolting 4788, Hanover, Germany           #
-- ########################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.atlas_core_package.all;

entity BOOT_MEM is
	port	(
				-- Host Interface --
				CLK_I           : in  std_logic; -- global clock line
				I_ADR_I         : in  std_logic_vector(15 downto 0); -- instruction adr
				I_EN_I          : in  std_logic; -- IR update
				I_DAT_O         : out std_logic_vector(15 downto 0); -- instruction out
				D_EN_I          : in  std_logic; -- access enable
				D_RW_I          : in  std_logic; -- read/write
				D_ADR_I         : in  std_logic_vector(15 downto 0); -- data adr
				D_DAT_I         : in  std_logic_vector(15 downto 0); -- data in
				D_DAT_O         : out std_logic_vector(15 downto 0)  -- data out
			);
end BOOT_MEM;

architecture BOOT_MEM_STRUCTURE of BOOT_MEM is

	-- Internal constants(configuration --
	constant mem_size_c      : natural := 2048; -- 2kB
	constant log2_mem_size_c : natural := log2(mem_size_c/2); -- address width (word boundary!)

	-- Memory Type --
	type mem_file_t is array (0 to (mem_size_c/2)-1) of std_logic_vector(15 downto 0); -- word mem!

	-- MEMORY IMAGE (Bootloader Program) --
	------------------------------------------------------
	constant BOOT_MEM_FILE_C : mem_file_t :=
    (
        000000 => x"bc0e", -- B
        000001 => x"bc04", -- B
        000002 => x"bc03", -- B
        000003 => x"bc02", -- B
        000004 => x"bc01", -- B
        000005 => x"c000", -- LDIL
        000006 => x"cc00", -- LDIH
        000007 => x"ec8a", -- MCR
        000008 => x"cc19", -- LDIH
        000009 => x"ed0f", -- MCR
        000010 => x"c52a", -- LDIL
        000011 => x"c907", -- LDIH
        000012 => x"be86", -- BL
        000013 => x"bc00", -- B
        000014 => x"ec11", -- MRC
        000015 => x"ec88", -- MCR
        000016 => x"ec8a", -- MCR
        000017 => x"c380", -- LDIL
        000018 => x"cff8", -- LDIH
        000019 => x"1c07", -- STSR
        000020 => x"2800", -- CLR
        000021 => x"ec08", -- MCR
        000022 => x"ec0b", -- MCR
        000023 => x"ec0e", -- MCR
        000024 => x"ec00", -- MRC
        000025 => x"ed88", -- MCR
        000026 => x"c002", -- LDIL
        000027 => x"ed8b", -- MCR
        000028 => x"c064", -- LDIL
        000029 => x"ed8d", -- MCR
        000030 => x"c901", -- LDIH
        000031 => x"ed2f", -- MCR
        000032 => x"ec17", -- MRC
        000033 => x"ec97", -- MRC
        000034 => x"c160", -- LDIL
        000035 => x"c909", -- LDIH
        000036 => x"c18f", -- LDIL
        000037 => x"0923", -- ADD
        000038 => x"29b3", -- CLR
        000039 => x"2a44", -- CLR
        000040 => x"100a", -- SUBS
        000041 => x"149b", -- SBCS
        000042 => x"9003", -- BMI
        000043 => x"0241", -- INC
        000044 => x"bdfc", -- B
        000045 => x"ed49", -- MCR
        000046 => x"ec22", -- MRC
        000047 => x"d406", -- SBR
        000048 => x"ed0a", -- MCR
        000049 => x"c538", -- LDIL
        000050 => x"c905", -- LDIH
        000051 => x"be5f", -- BL
        000052 => x"c12e", -- LDIL
        000053 => x"c906", -- LDIH
        000054 => x"be5c", -- BL
        000055 => x"ee11", -- MRC
        000056 => x"be5e", -- BL
        000057 => x"c13e", -- LDIL
        000058 => x"c906", -- LDIH
        000059 => x"be57", -- BL
        000060 => x"ee97", -- MRC
        000061 => x"ee17", -- MRC
        000062 => x"be58", -- BL
        000063 => x"0250", -- MOV
        000064 => x"be56", -- BL
        000065 => x"be52", -- BL
        000066 => x"ec27", -- MRC
        000067 => x"c083", -- LDIL
        000068 => x"2001", -- AND
        000069 => x"c330", -- LDIL
        000070 => x"0b60", -- ADD
        000071 => x"bc0f", -- B
        000072 => x"c55e", -- LDIL
        000073 => x"c906", -- LDIH
        000074 => x"be48", -- BL
        000075 => x"c14e", -- LDIL
        000076 => x"c907", -- LDIH
        000077 => x"be45", -- BL
        000078 => x"c514", -- LDIL
        000079 => x"c907", -- LDIH
        000080 => x"be42", -- BL
        000081 => x"be44", -- BL
        000082 => x"0300", -- MOV
        000083 => x"0080", -- MOV
        000084 => x"be40", -- BL
        000085 => x"be3e", -- BL
        000086 => x"c0b0", -- LDIL
        000087 => x"181e", -- CMP
        000088 => x"81f0", -- BEQ
        000089 => x"c0b1", -- LDIL
        000090 => x"181e", -- CMP
        000091 => x"809b", -- BEQ
        000092 => x"c0b2", -- LDIL
        000093 => x"181e", -- CMP
        000094 => x"8064", -- BEQ
        000095 => x"c0b3", -- LDIL
        000096 => x"181e", -- CMP
        000097 => x"802b", -- BEQ
        000098 => x"c0b4", -- LDIL
        000099 => x"181e", -- CMP
        000100 => x"8033", -- BEQ
        000101 => x"c0bf", -- LDIL
        000102 => x"181e", -- CMP
        000103 => x"8405", -- BNE
        000104 => x"c102", -- LDIL
        000105 => x"c901", -- LDIH
        000106 => x"be28", -- BL
        000107 => x"bde3", -- B
        000108 => x"c2be", -- LDIL
        000109 => x"ca83", -- LDIH
        000110 => x"c0f0", -- LDIL
        000111 => x"181e", -- CMP
        000112 => x"f705", -- RBAEQ
        000113 => x"c0e4", -- LDIL
        000114 => x"181e", -- CMP
        000115 => x"80f1", -- BEQ
        000116 => x"c2e4", -- LDIL
        000117 => x"ca85", -- LDIH
        000118 => x"c0f7", -- LDIL
        000119 => x"181e", -- CMP
        000120 => x"f705", -- RBAEQ
        000121 => x"c0f2", -- LDIL
        000122 => x"181e", -- CMP
        000123 => x"85d3", -- BNE
        000124 => x"2800", -- CLR
        000125 => x"c080", -- LDIL
        000126 => x"cc80", -- LDIH
        000127 => x"ec99", -- MCR
        000128 => x"3400", -- GT
        000129 => x"4b65", -- .DW
        000130 => x"6570", -- .DW
        000131 => x"696e", -- .DW
        000132 => x"2720", -- .DW
        000133 => x"6974", -- .DW
        000134 => x"2063", -- .DW
        000135 => x"6f75", -- .DW
        000136 => x"6e74", -- .DW
        000137 => x"7279", -- .DW
        000138 => x"210d", -- .DW
        000139 => x"0a00", -- .DW
        000140 => x"c14e", -- LDIL
        000141 => x"c906", -- LDIH
        000142 => x"be04", -- BL
        000143 => x"2800", -- CLR
        000144 => x"2100", -- STUB
        000145 => x"bca7", -- B
        000146 => x"bc9c", -- B
        000147 => x"bc9c", -- B
        000148 => x"bc9c", -- B
        000149 => x"bc9c", -- B
        000150 => x"bc9f", -- B
        000151 => x"c52e", -- LDIL
        000152 => x"c906", -- LDIH
        000153 => x"be95", -- BL
        000154 => x"be9d", -- BL
        000155 => x"edca", -- MCR
        000156 => x"be9b", -- BL
        000157 => x"edc9", -- MCR
        000158 => x"c426", -- LDIL
        000159 => x"c805", -- LDIH
        000160 => x"3404", -- GTL
        000161 => x"be8e", -- BL
        000162 => x"be94", -- BL
        000163 => x"c47e", -- LDIL
        000164 => x"cc4a", -- LDIH
        000165 => x"180e", -- CMP
        000166 => x"848d", -- BNE
        000167 => x"be8f", -- BL
        000168 => x"3f64", -- SFT
        000169 => x"2066", -- STUB
        000170 => x"be8c", -- BL
        000171 => x"20e6", -- STUB
        000172 => x"be8a", -- BL
        000173 => x"2166", -- STUB
        000174 => x"be88", -- BL
        000175 => x"21e6", -- STUB
        000176 => x"be86", -- BL
        000177 => x"2266", -- STUB
        000178 => x"be84", -- BL
        000179 => x"22e6", -- STUB
        000180 => x"be82", -- BL
        000181 => x"2366", -- STUB
        000182 => x"c280", -- LDIL
        000183 => x"ecda", -- MCR
        000184 => x"ec5d", -- MCR
        000185 => x"be7d", -- BL
        000186 => x"7f5a", -- STR
        000187 => x"ec05", -- MRC
        000188 => x"2806", -- EOR
        000189 => x"ec0d", -- MCR
        000190 => x"2400", -- LDUB
        000191 => x"1858", -- CMP
        000192 => x"85f9", -- BNE
        000193 => x"bc5a", -- B
        000194 => x"c14e", -- LDIL
        000195 => x"c906", -- LDIH
        000196 => x"be6a", -- BL
        000197 => x"c100", -- LDIL
        000198 => x"be29", -- BL
        000199 => x"c47e", -- LDIL
        000200 => x"cc4a", -- LDIH
        000201 => x"180d", -- CMP
        000202 => x"8469", -- BNE
        000203 => x"c102", -- LDIL
        000204 => x"be23", -- BL
        000205 => x"3ed4", -- SFT
        000206 => x"2055", -- STUB
        000207 => x"c104", -- LDIL
        000208 => x"be1f", -- BL
        000209 => x"20d5", -- STUB
        000210 => x"c106", -- LDIL
        000211 => x"be1c", -- BL
        000212 => x"2155", -- STUB
        000213 => x"c108", -- LDIL
        000214 => x"be19", -- BL
        000215 => x"21d5", -- STUB
        000216 => x"c10a", -- LDIL
        000217 => x"be16", -- BL
        000218 => x"2255", -- STUB
        000219 => x"c10c", -- LDIL
        000220 => x"be13", -- BL
        000221 => x"22d5", -- STUB
        000222 => x"c10e", -- LDIL
        000223 => x"be10", -- BL
        000224 => x"2355", -- STUB
        000225 => x"c200", -- LDIL
        000226 => x"ecca", -- MCR
        000227 => x"ec4d", -- MCR
        000228 => x"c010", -- LDIL
        000229 => x"0940", -- ADD
        000230 => x"be09", -- BL
        000231 => x"7eca", -- STR
        000232 => x"ec05", -- MRC
        000233 => x"2805", -- EOR
        000234 => x"ec0d", -- MCR
        000235 => x"2400", -- LDUB
        000236 => x"1848", -- CMP
        000237 => x"85f7", -- BNE
        000238 => x"bc2d", -- B
        000239 => x"0370", -- MOV
        000240 => x"be42", -- BL
        000241 => x"3eb0", -- SFT
        000242 => x"0121", -- INC
        000243 => x"be3f", -- BL
        000244 => x"26d3", -- ORR
        000245 => x"3460", -- RET
        000246 => x"c166", -- LDIL
        000247 => x"c906", -- LDIH
        000248 => x"be36", -- BL
        000249 => x"be38", -- BL
        000250 => x"3c80", -- SFT
        000251 => x"be36", -- BL
        000252 => x"2490", -- ORR
        000253 => x"c47e", -- LDIL
        000254 => x"cc4a", -- LDIH
        000255 => x"1818", -- CMP
        000256 => x"8433", -- BNE
        000257 => x"be27", -- BL
        000258 => x"3c94", -- SFT
        000259 => x"2011", -- STUB
        000260 => x"be24", -- BL
        000261 => x"2091", -- STUB
        000262 => x"be22", -- BL
        000263 => x"2111", -- STUB
        000264 => x"be20", -- BL
        000265 => x"2191", -- STUB
        000266 => x"be1e", -- BL
        000267 => x"2211", -- STUB
        000268 => x"be1c", -- BL
        000269 => x"2291", -- STUB
        000270 => x"be1a", -- BL
        000271 => x"2311", -- STUB
        000272 => x"2ad5", -- CLR
        000273 => x"ecda", -- MCR
        000274 => x"ec5d", -- MCR
        000275 => x"be15", -- BL
        000276 => x"7cda", -- STR
        000277 => x"ec05", -- MRC
        000278 => x"2801", -- EOR
        000279 => x"ec0d", -- MCR
        000280 => x"2400", -- LDUB
        000281 => x"1858", -- CMP
        000282 => x"85f9", -- BNE
        000283 => x"ec11", -- MRC
        000284 => x"ec8a", -- MCR
        000285 => x"c50c", -- LDIL
        000286 => x"c906", -- LDIH
        000287 => x"be0f", -- BL
        000288 => x"ec05", -- MRC
        000289 => x"2491", -- LDUB
        000290 => x"1809", -- CMP
        000291 => x"8015", -- BEQ
        000292 => x"c538", -- LDIL
        000293 => x"c907", -- LDIH
        000294 => x"be08", -- BL
        000295 => x"bccb", -- B
        000296 => x"0370", -- MOV
        000297 => x"be08", -- BL
        000298 => x"3c80", -- SFT
        000299 => x"be06", -- BL
        000300 => x"2490", -- ORR
        000301 => x"3460", -- RET
        000302 => x"bcc7", -- B
        000303 => x"bcd0", -- B
        000304 => x"bcd4", -- B
        000305 => x"bcd8", -- B
        000306 => x"bc6b", -- B
        000307 => x"bcbc", -- B
        000308 => x"bd1a", -- B
        000309 => x"bc69", -- B
        000310 => x"bcbe", -- B
        000311 => x"bcd7", -- B
        000312 => x"c54c", -- LDIL
        000313 => x"c906", -- LDIH
        000314 => x"bebb", -- BL
        000315 => x"ee05", -- MRC
        000316 => x"bef7", -- BL
        000317 => x"bec2", -- BL
        000318 => x"c17c", -- LDIL
        000319 => x"c906", -- LDIH
        000320 => x"beb5", -- BL
        000321 => x"24aa", -- LDUBS
        000322 => x"8010", -- BEQ
        000323 => x"c0a2", -- LDIL
        000324 => x"bec0", -- BL
        000325 => x"24a2", -- LDUB
        000326 => x"be18", -- BL
        000327 => x"24b3", -- LDUB
        000328 => x"be16", -- BL
        000329 => x"24c4", -- LDUB
        000330 => x"be14", -- BL
        000331 => x"24d5", -- LDUB
        000332 => x"be12", -- BL
        000333 => x"24e6", -- LDUB
        000334 => x"be10", -- BL
        000335 => x"c0a2", -- LDIL
        000336 => x"beb4", -- BL
        000337 => x"beae", -- BL
        000338 => x"bead", -- BL
        000339 => x"c080", -- LDIL
        000340 => x"ccc0", -- LDIH
        000341 => x"1c01", -- STSR
        000342 => x"2800", -- CLR
        000343 => x"ed0f", -- MCR
        000344 => x"ec88", -- MCR
        000345 => x"ec8b", -- MCR
        000346 => x"ec8c", -- MCR
        000347 => x"ec8a", -- MCR
        000348 => x"ec89", -- MCR
        000349 => x"3400", -- GT
        000350 => x"0370", -- MOV
        000351 => x"3c90", -- SFT
        000352 => x"bea4", -- BL
        000353 => x"3c90", -- SFT
        000354 => x"bea2", -- BL
        000355 => x"3460", -- RET
        000356 => x"c520", -- LDIL
        000357 => x"c906", -- LDIH
        000358 => x"be8f", -- BL
        000359 => x"bea7", -- BL
        000360 => x"c526", -- LDIL
        000361 => x"c905", -- LDIH
        000362 => x"3424", -- GTL
        000363 => x"ecca", -- MCR
        000364 => x"be93", -- BL
        000365 => x"c280", -- LDIL
        000366 => x"c00f", -- LDIL
        000367 => x"2058", -- ANDS
        000368 => x"840a", -- BNE
        000369 => x"be8e", -- BL
        000370 => x"c0a4", -- LDIL
        000371 => x"be91", -- BL
        000372 => x"0250", -- MOV
        000373 => x"bebe", -- BL
        000374 => x"c0ba", -- LDIL
        000375 => x"be8d", -- BL
        000376 => x"c0a0", -- LDIL
        000377 => x"be8b", -- BL
        000378 => x"7a5a", -- LDR
        000379 => x"c0a0", -- LDIL
        000380 => x"be88", -- BL
        000381 => x"beb6", -- BL
        000382 => x"c00f", -- LDIL
        000383 => x"2058", -- ANDS
        000384 => x"8414", -- BNE
        000385 => x"c0a0", -- LDIL
        000386 => x"be82", -- BL
        000387 => x"be81", -- BL
        000388 => x"c010", -- LDIL
        000389 => x"1250", -- SUB
        000390 => x"c470", -- LDIL
        000391 => x"2240", -- AND
        000392 => x"78c9", -- LDR
        000393 => x"3c90", -- SFT
        000394 => x"c880", -- LDIH
        000395 => x"c020", -- LDIL
        000396 => x"1818", -- CMP
        000397 => x"a402", -- BLS
        000398 => x"c0ae", -- LDIL
        000399 => x"be75", -- BL
        000400 => x"c08f", -- LDIL
        000401 => x"2014", -- AND
        000402 => x"3409", -- TEQ
        000403 => x"85f5", -- BNE
        000404 => x"ec20", -- MRC
        000405 => x"dc0f", -- STB
        000406 => x"b804", -- BTS
        000407 => x"c5fe", -- LDIL
        000408 => x"343d", -- TEQ
        000409 => x"85d5", -- BNE
        000410 => x"be6f", -- BL
        000411 => x"2800", -- CLR
        000412 => x"3400", -- GT
        000413 => x"bc56", -- B
        000414 => x"bc95", -- B
        000415 => x"c001", -- LDIL
        000416 => x"ed0c", -- MCR
        000417 => x"c050", -- LDIL
        000418 => x"c83f", -- LDIH
        000419 => x"ed0a", -- MCR
        000420 => x"c000", -- LDIL
        000421 => x"c801", -- LDIH
        000422 => x"beab", -- BL
        000423 => x"c158", -- LDIL
        000424 => x"c906", -- LDIH
        000425 => x"be4c", -- BL
        000426 => x"c166", -- LDIL
        000427 => x"c906", -- LDIH
        000428 => x"be49", -- BL
        000429 => x"be5c", -- BL
        000430 => x"3c80", -- SFT
        000431 => x"be5a", -- BL
        000432 => x"2410", -- ORR
        000433 => x"c4fe", -- LDIL
        000434 => x"ccca", -- LDIH
        000435 => x"1809", -- CMP
        000436 => x"843b", -- BNE
        000437 => x"c100", -- LDIL
        000438 => x"c6fe", -- LDIL
        000439 => x"ceca", -- LDIH
        000440 => x"be30", -- BL
        000441 => x"be50", -- BL
        000442 => x"3c80", -- SFT
        000443 => x"be4e", -- BL
        000444 => x"2690", -- ORR
        000445 => x"3ed4", -- SFT
        000446 => x"2055", -- STUB
        000447 => x"c102", -- LDIL
        000448 => x"be28", -- BL
        000449 => x"be48", -- BL
        000450 => x"3c80", -- SFT
        000451 => x"be46", -- BL
        000452 => x"2690", -- ORR
        000453 => x"20d5", -- STUB
        000454 => x"c104", -- LDIL
        000455 => x"be21", -- BL
        000456 => x"c106", -- LDIL
        000457 => x"be40", -- BL
        000458 => x"0180", -- MOV
        000459 => x"be8c", -- BL
        000460 => x"0121", -- INC
        000461 => x"c010", -- LDIL
        000462 => x"1828", -- CMP
        000463 => x"85fa", -- BNE
        000464 => x"c110", -- LDIL
        000465 => x"2ad5", -- CLR
        000466 => x"be37", -- BL
        000467 => x"0180", -- MOV
        000468 => x"be83", -- BL
        000469 => x"0121", -- INC
        000470 => x"2400", -- LDUB
        000471 => x"02d1", -- INC
        000472 => x"1858", -- CMP
        000473 => x"85f9", -- BNE
        000474 => x"c001", -- LDIL
        000475 => x"ed0c", -- MCR
        000476 => x"c050", -- LDIL
        000477 => x"c83f", -- LDIH
        000478 => x"ed0a", -- MCR
        000479 => x"c00c", -- LDIL
        000480 => x"c801", -- LDIH
        000481 => x"be70", -- BL
        000482 => x"c50c", -- LDIL
        000483 => x"c906", -- LDIH
        000484 => x"be11", -- BL
        000485 => x"c690", -- LDIL
        000486 => x"ca80", -- LDIH
        000487 => x"3450", -- GT
        000488 => x"0370", -- MOV
        000489 => x"3dd0", -- SFT
        000490 => x"be6d", -- BL
        000491 => x"0121", -- INC
        000492 => x"01d0", -- MOV
        000493 => x"be6a", -- BL
        000494 => x"3460", -- RET
        000495 => x"c51c", -- LDIL
        000496 => x"c907", -- LDIH
        000497 => x"be04", -- BL
        000498 => x"bcba", -- B
        000499 => x"bc94", -- B
        000500 => x"bca5", -- B
        000501 => x"01f0", -- MOV
        000502 => x"7829", -- LDR
        000503 => x"c080", -- LDIL
        000504 => x"ccff", -- LDIH
        000505 => x"2081", -- AND
        000506 => x"3c98", -- SFTS
        000507 => x"8003", -- BEQ
        000508 => x"be08", -- BL
        000509 => x"bdf9", -- B
        000510 => x"3430", -- RET
        000511 => x"0170", -- MOV
        000512 => x"c08d", -- LDIL
        000513 => x"be03", -- BL
        000514 => x"c08a", -- LDIL
        000515 => x"03a0", -- MOV
        000516 => x"ec22", -- MRC
        000517 => x"dc05", -- STB
        000518 => x"b9fe", -- BTS
        000519 => x"ed18", -- MCR
        000520 => x"3470", -- RET
        000521 => x"ec20", -- MRC
        000522 => x"dc8f", -- STBI
        000523 => x"b9fe", -- BTS
        000524 => x"c800", -- LDIH
        000525 => x"3470", -- RET
        000526 => x"0170", -- MOV
        000527 => x"c200", -- LDIL
        000528 => x"c184", -- LDIL
        000529 => x"bff8", -- BL
        000530 => x"c0c6", -- LDIL
        000531 => x"1809", -- CMP
        000532 => x"9003", -- BMI
        000533 => x"c0a0", -- LDIL
        000534 => x"1001", -- SUB
        000535 => x"c0b0", -- LDIL
        000536 => x"1809", -- CMP
        000537 => x"91f8", -- BMI
        000538 => x"c0c6", -- LDIL
        000539 => x"1818", -- CMP
        000540 => x"91f5", -- BMI
        000541 => x"c0b9", -- LDIL
        000542 => x"1818", -- CMP
        000543 => x"a404", -- BLS
        000544 => x"c0c1", -- LDIL
        000545 => x"1809", -- CMP
        000546 => x"a1ef", -- BHI
        000547 => x"0080", -- MOV
        000548 => x"bfe0", -- BL
        000549 => x"c030", -- LDIL
        000550 => x"1090", -- SUB
        000551 => x"c009", -- LDIL
        000552 => x"1809", -- CMP
        000553 => x"a402", -- BLS
        000554 => x"0497", -- DEC
        000555 => x"3e42", -- SFT
        000556 => x"3e42", -- SFT
        000557 => x"3e42", -- SFT
        000558 => x"3e42", -- SFT
        000559 => x"2641", -- ORR
        000560 => x"05b9", -- DECS
        000561 => x"85e0", -- BNE
        000562 => x"3420", -- RET
        000563 => x"0370", -- MOV
        000564 => x"3d42", -- SFT
        000565 => x"3d22", -- SFT
        000566 => x"3d22", -- SFT
        000567 => x"3d22", -- SFT
        000568 => x"be0f", -- BL
        000569 => x"bfcb", -- BL
        000570 => x"3d40", -- SFT
        000571 => x"be0c", -- BL
        000572 => x"bfc8", -- BL
        000573 => x"3d45", -- SFT
        000574 => x"3d25", -- SFT
        000575 => x"3d25", -- SFT
        000576 => x"3d25", -- SFT
        000577 => x"be06", -- BL
        000578 => x"bfc2", -- BL
        000579 => x"0140", -- MOV
        000580 => x"be03", -- BL
        000581 => x"bfbf", -- BL
        000582 => x"3460", -- RET
        000583 => x"c08f", -- LDIL
        000584 => x"2121", -- AND
        000585 => x"c089", -- LDIL
        000586 => x"181a", -- CMP
        000587 => x"8803", -- BCS
        000588 => x"c0b0", -- LDIL
        000589 => x"bc02", -- B
        000590 => x"c0b7", -- LDIL
        000591 => x"0892", -- ADD
        000592 => x"3470", -- RET
        000593 => x"ed0b", -- MCR
        000594 => x"ec22", -- MRC
        000595 => x"dc03", -- STB
        000596 => x"b9fe", -- BTS
        000597 => x"ec23", -- MRC
        000598 => x"3470", -- RET
        000599 => x"00f0", -- MOV
        000600 => x"c050", -- LDIL
        000601 => x"c837", -- LDIH
        000602 => x"ed0a", -- MCR
        000603 => x"c001", -- LDIL
        000604 => x"ed0c", -- MCR
        000605 => x"c006", -- LDIL
        000606 => x"bff3", -- BL
        000607 => x"c050", -- LDIL
        000608 => x"c83f", -- LDIH
        000609 => x"ed0a", -- MCR
        000610 => x"c000", -- LDIL
        000611 => x"c805", -- LDIH
        000612 => x"bfed", -- BL
        000613 => x"dc01", -- STB
        000614 => x"b805", -- BTS
        000615 => x"c548", -- LDIL
        000616 => x"c907", -- LDIH
        000617 => x"bf8c", -- BL
        000618 => x"bc42", -- B
        000619 => x"c040", -- LDIL
        000620 => x"c83f", -- LDIH
        000621 => x"ed0a", -- MCR
        000622 => x"c001", -- LDIL
        000623 => x"ed0c", -- MCR
        000624 => x"3c20", -- SFT
        000625 => x"c802", -- LDIH
        000626 => x"bfdf", -- BL
        000627 => x"03a0", -- MOV
        000628 => x"cb80", -- LDIH
        000629 => x"3ff0", -- SFT
        000630 => x"0030", -- MOV
        000631 => x"c800", -- LDIH
        000632 => x"2407", -- ORR
        000633 => x"bfd8", -- BL
        000634 => x"2800", -- CLR
        000635 => x"ed0c", -- MCR
        000636 => x"c050", -- LDIL
        000637 => x"c83f", -- LDIH
        000638 => x"ed0a", -- MCR
        000639 => x"c001", -- LDIL
        000640 => x"ed0c", -- MCR
        000641 => x"c000", -- LDIL
        000642 => x"c805", -- LDIH
        000643 => x"bfce", -- BL
        000644 => x"dc00", -- STB
        000645 => x"b9fc", -- BTS
        000646 => x"3410", -- RET
        000647 => x"00f0", -- MOV
        000648 => x"c040", -- LDIL
        000649 => x"c83f", -- LDIH
        000650 => x"ed0a", -- MCR
        000651 => x"c001", -- LDIL
        000652 => x"ed0c", -- MCR
        000653 => x"3c20", -- SFT
        000654 => x"c803", -- LDIH
        000655 => x"bfc2", -- BL
        000656 => x"0020", -- MOV
        000657 => x"c800", -- LDIH
        000658 => x"3c00", -- SFT
        000659 => x"bfbe", -- BL
        000660 => x"29b3", -- CLR
        000661 => x"ed3c", -- MCR
        000662 => x"0180", -- MOV
        000663 => x"c980", -- LDIH
        000664 => x"3410", -- RET
        000665 => x"e5b0", -- CDP
        000666 => x"ec30", -- MRC
        000667 => x"dc06", -- STB
        000668 => x"b9fe", -- BTS
        000669 => x"c306", -- LDIL
        000670 => x"200e", -- ANDS
        000671 => x"840a", -- BNE
        000672 => x"ecb1", -- MRC
        000673 => x"ef32", -- MRC
        000674 => x"2800", -- CLR
        000675 => x"009a", -- INCS
        000676 => x"0f60", -- ADC
        000677 => x"ed99", -- MCR
        000678 => x"edea", -- MCR
        000679 => x"ef34", -- MRC
        000680 => x"3470", -- RET
        000681 => x"c55a", -- LDIL
        000682 => x"c907", -- LDIH
        000683 => x"bf4a", -- BL
        000684 => x"c568", -- LDIL
        000685 => x"c907", -- LDIH
        000686 => x"bf47", -- BL
        000687 => x"bf5a", -- BL
        000688 => x"2800", -- CLR
        000689 => x"3400", -- GT
        000690 => x"c52e", -- LDIL
        000691 => x"c906", -- LDIH
        000692 => x"bf41", -- BL
        000693 => x"bf59", -- BL
        000694 => x"edca", -- MCR
        000695 => x"bf57", -- BL
        000696 => x"edc9", -- MCR
        000697 => x"be1a", -- BL
        000698 => x"bf45", -- BL
        000699 => x"c53c", -- LDIL
        000700 => x"c906", -- LDIH
        000701 => x"bf38", -- BL
        000702 => x"bf50", -- BL
        000703 => x"02c0", -- MOV
        000704 => x"be13", -- BL
        000705 => x"345d", -- TEQ
        000706 => x"800d", -- BEQ
        000707 => x"06d1", -- DEC
        000708 => x"bf3b", -- BL
        000709 => x"bfd4", -- BL
        000710 => x"c558", -- LDIL
        000711 => x"c906", -- LDIH
        000712 => x"bf2d", -- BL
        000713 => x"0260", -- MOV
        000714 => x"bf69", -- BL
        000715 => x"eca0", -- MRC
        000716 => x"dc1f", -- STB
        000717 => x"b802", -- BTS
        000718 => x"bdf3", -- B
        000719 => x"bf30", -- BL
        000720 => x"c69c", -- LDIL
        000721 => x"ca80", -- LDIH
        000722 => x"3450", -- GT
        000723 => x"0170", -- MOV
        000724 => x"bf35", -- BL
        000725 => x"c08d", -- LDIL
        000726 => x"1809", -- CMP
        000727 => x"f702", -- RBAEQ
        000728 => x"c088", -- LDIL
        000729 => x"1809", -- CMP
        000730 => x"81f5", -- BEQ
        000731 => x"bdf9", -- B
        000732 => x"0d0a", -- .DW
        000733 => x"0d0a", -- .DW
        000734 => x"4174", -- .DW
        000735 => x"6c61", -- .DW
        000736 => x"732d", -- .DW
        000737 => x"324b", -- .DW
        000738 => x"2042", -- .DW
        000739 => x"6f6f", -- .DW
        000740 => x"746c", -- .DW
        000741 => x"6f61", -- .DW
        000742 => x"6465", -- .DW
        000743 => x"7220", -- .DW
        000744 => x"2d20", -- .DW
        000745 => x"5632", -- .DW
        000746 => x"3031", -- .DW
        000747 => x"3430", -- .DW
        000748 => x"3431", -- .DW
        000749 => x"340d", -- .DW
        000750 => x"0a62", -- .DW
        000751 => x"7920", -- .DW
        000752 => x"5374", -- .DW
        000753 => x"6570", -- .DW
        000754 => x"6861", -- .DW
        000755 => x"6e20", -- .DW
        000756 => x"4e6f", -- .DW
        000757 => x"6c74", -- .DW
        000758 => x"696e", -- .DW
        000759 => x"672c", -- .DW
        000760 => x"2073", -- .DW
        000761 => x"746e", -- .DW
        000762 => x"6f6c", -- .DW
        000763 => x"7469", -- .DW
        000764 => x"6e67", -- .DW
        000765 => x"4067", -- .DW
        000766 => x"6d61", -- .DW
        000767 => x"696c", -- .DW
        000768 => x"2e63", -- .DW
        000769 => x"6f6d", -- .DW
        000770 => x"0d0a", -- .DW
        000771 => x"7777", -- .DW
        000772 => x"772e", -- .DW
        000773 => x"6f70", -- .DW
        000774 => x"656e", -- .DW
        000775 => x"636f", -- .DW
        000776 => x"7265", -- .DW
        000777 => x"732e", -- .DW
        000778 => x"6f72", -- .DW
        000779 => x"672f", -- .DW
        000780 => x"7072", -- .DW
        000781 => x"6f6a", -- .DW
        000782 => x"6563", -- .DW
        000783 => x"742c", -- .DW
        000784 => x"6174", -- .DW
        000785 => x"6c61", -- .DW
        000786 => x"735f", -- .DW
        000787 => x"636f", -- .DW
        000788 => x"7265", -- .DW
        000789 => x"0d0a", -- .DW
        000790 => x"0000", -- .DW
        000791 => x"0d0a", -- .DW
        000792 => x"426f", -- .DW
        000793 => x"6f74", -- .DW
        000794 => x"2070", -- .DW
        000795 => x"6167", -- .DW
        000796 => x"653a", -- .DW
        000797 => x"2030", -- .DW
        000798 => x"7800", -- .DW
        000799 => x"0d0a", -- .DW
        000800 => x"436c", -- .DW
        000801 => x"6f63", -- .DW
        000802 => x"6b28", -- .DW
        000803 => x"487a", -- .DW
        000804 => x"293a", -- .DW
        000805 => x"2030", -- .DW
        000806 => x"7800", -- .DW
        000807 => x"426f", -- .DW
        000808 => x"6f74", -- .DW
        000809 => x"696e", -- .DW
        000810 => x"670d", -- .DW
        000811 => x"0a00", -- .DW
        000812 => x"4275", -- .DW
        000813 => x"726e", -- .DW
        000814 => x"2045", -- .DW
        000815 => x"4550", -- .DW
        000816 => x"524f", -- .DW
        000817 => x"4d0d", -- .DW
        000818 => x"0a00", -- .DW
        000819 => x"5761", -- .DW
        000820 => x"6974", -- .DW
        000821 => x"696e", -- .DW
        000822 => x"6720", -- .DW
        000823 => x"666f", -- .DW
        000824 => x"7220", -- .DW
        000825 => x"6461", -- .DW
        000826 => x"7461", -- .DW
        000827 => x"2e2e", -- .DW
        000828 => x"2e0d", -- .DW
        000829 => x"0a00", -- .DW
        000830 => x"5374", -- .DW
        000831 => x"6172", -- .DW
        000832 => x"7469", -- .DW
        000833 => x"6e67", -- .DW
        000834 => x"2069", -- .DW
        000835 => x"6d61", -- .DW
        000836 => x"6765", -- .DW
        000837 => x"2000", -- .DW
        000838 => x"446f", -- .DW
        000839 => x"776e", -- .DW
        000840 => x"6c6f", -- .DW
        000841 => x"6164", -- .DW
        000842 => x"2063", -- .DW
        000843 => x"6f6d", -- .DW
        000844 => x"706c", -- .DW
        000845 => x"6574", -- .DW
        000846 => x"650d", -- .DW
        000847 => x"0a00", -- .DW
        000848 => x"5061", -- .DW
        000849 => x"6765", -- .DW
        000850 => x"2028", -- .DW
        000851 => x"3468", -- .DW
        000852 => x"293a", -- .DW
        000853 => x"2024", -- .DW
        000854 => x"0000", -- .DW
        000855 => x"4164", -- .DW
        000856 => x"6472", -- .DW
        000857 => x"2028", -- .DW
        000858 => x"3868", -- .DW
        000859 => x"293a", -- .DW
        000860 => x"2024", -- .DW
        000861 => x"0000", -- .DW
        000862 => x"2377", -- .DW
        000863 => x"6f72", -- .DW
        000864 => x"6473", -- .DW
        000865 => x"2028", -- .DW
        000866 => x"3468", -- .DW
        000867 => x"293a", -- .DW
        000868 => x"2024", -- .DW
        000869 => x"0000", -- .DW
        000870 => x"4368", -- .DW
        000871 => x"6563", -- .DW
        000872 => x"6b73", -- .DW
        000873 => x"756d", -- .DW
        000874 => x"3a20", -- .DW
        000875 => x"2400", -- .DW
        000876 => x"202d", -- .DW
        000877 => x"3e20", -- .DW
        000878 => x"2400", -- .DW
        000879 => x"0d0a", -- .DW
        000880 => x"636d", -- .DW
        000881 => x"642f", -- .DW
        000882 => x"626f", -- .DW
        000883 => x"6f74", -- .DW
        000884 => x"2d73", -- .DW
        000885 => x"7769", -- .DW
        000886 => x"7463", -- .DW
        000887 => x"683a", -- .DW
        000888 => x"0d0a", -- .DW
        000889 => x"2030", -- .DW
        000890 => x"2f27", -- .DW
        000891 => x"3030", -- .DW
        000892 => x"273a", -- .DW
        000893 => x"2052", -- .DW
        000894 => x"6573", -- .DW
        000895 => x"7461", -- .DW
        000896 => x"7274", -- .DW
        000897 => x"2063", -- .DW
        000898 => x"6f6e", -- .DW
        000899 => x"736f", -- .DW
        000900 => x"6c65", -- .DW
        000901 => x"0d0a", -- .DW
        000902 => x"2031", -- .DW
        000903 => x"2f27", -- .DW
        000904 => x"3031", -- .DW
        000905 => x"273a", -- .DW
        000906 => x"2042", -- .DW
        000907 => x"6f6f", -- .DW
        000908 => x"7420", -- .DW
        000909 => x"5541", -- .DW
        000910 => x"5254", -- .DW
        000911 => x"0d0a", -- .DW
        000912 => x"2032", -- .DW
        000913 => x"2f27", -- .DW
        000914 => x"3130", -- .DW
        000915 => x"273a", -- .DW
        000916 => x"2042", -- .DW
        000917 => x"6f6f", -- .DW
        000918 => x"7420", -- .DW
        000919 => x"4545", -- .DW
        000920 => x"5052", -- .DW
        000921 => x"4f4d", -- .DW
        000922 => x"0d0a", -- .DW
        000923 => x"2033", -- .DW
        000924 => x"2f27", -- .DW
        000925 => x"3131", -- .DW
        000926 => x"273a", -- .DW
        000927 => x"2042", -- .DW
        000928 => x"6f6f", -- .DW
        000929 => x"7420", -- .DW
        000930 => x"6d65", -- .DW
        000931 => x"6d6f", -- .DW
        000932 => x"7279", -- .DW
        000933 => x"0d0a", -- .DW
        000934 => x"0000", -- .DW
        000935 => x"2034", -- .DW
        000936 => x"3a20", -- .DW
        000937 => x"426f", -- .DW
        000938 => x"6f74", -- .DW
        000939 => x"2057", -- .DW
        000940 => x"420d", -- .DW
        000941 => x"0a20", -- .DW
        000942 => x"703a", -- .DW
        000943 => x"2042", -- .DW
        000944 => x"7572", -- .DW
        000945 => x"6e20", -- .DW
        000946 => x"4545", -- .DW
        000947 => x"5052", -- .DW
        000948 => x"4f4d", -- .DW
        000949 => x"0d0a", -- .DW
        000950 => x"2064", -- .DW
        000951 => x"3a20", -- .DW
        000952 => x"5241", -- .DW
        000953 => x"4d20", -- .DW
        000954 => x"6475", -- .DW
        000955 => x"6d70", -- .DW
        000956 => x"0d0a", -- .DW
        000957 => x"2072", -- .DW
        000958 => x"3a20", -- .DW
        000959 => x"5265", -- .DW
        000960 => x"7365", -- .DW
        000961 => x"740d", -- .DW
        000962 => x"0a20", -- .DW
        000963 => x"773a", -- .DW
        000964 => x"2057", -- .DW
        000965 => x"4220", -- .DW
        000966 => x"6475", -- .DW
        000967 => x"6d70", -- .DW
        000968 => x"0d0a", -- .DW
        000969 => x"0000", -- .DW
        000970 => x"636d", -- .DW
        000971 => x"643a", -- .DW
        000972 => x"3e20", -- .DW
        000973 => x"0000", -- .DW
        000974 => x"494d", -- .DW
        000975 => x"4147", -- .DW
        000976 => x"4520", -- .DW
        000977 => x"4552", -- .DW
        000978 => x"5221", -- .DW
        000979 => x"0d0a", -- .DW
        000980 => x"0000", -- .DW
        000981 => x"0d0a", -- .DW
        000982 => x"4952", -- .DW
        000983 => x"5120", -- .DW
        000984 => x"4552", -- .DW
        000985 => x"5221", -- .DW
        000986 => x"0d0a", -- .DW
        000987 => x"0000", -- .DW
        000988 => x"4348", -- .DW
        000989 => x"4543", -- .DW
        000990 => x"4b53", -- .DW
        000991 => x"554d", -- .DW
        000992 => x"2045", -- .DW
        000993 => x"5252", -- .DW
        000994 => x"210d", -- .DW
        000995 => x"0a00", -- .DW
        000996 => x"5350", -- .DW
        000997 => x"492f", -- .DW
        000998 => x"4545", -- .DW
        000999 => x"5052", -- .DW
        001000 => x"4f4d", -- .DW
        001001 => x"2045", -- .DW
        001002 => x"5252", -- .DW
        001003 => x"210d", -- .DW
        001004 => x"0a00", -- .DW
        001005 => x"5742", -- .DW
        001006 => x"2042", -- .DW
        001007 => x"5553", -- .DW
        001008 => x"2045", -- .DW
        001009 => x"5252", -- .DW
        001010 => x"210d", -- .DW
        001011 => x"0a00", -- .DW
        001012 => x"5072", -- .DW
        001013 => x"6573", -- .DW
        001014 => x"7320", -- .DW
        001015 => x"616e", -- .DW
        001016 => x"7920", -- .DW
        001017 => x"6b65", -- .DW
        001018 => x"790d", -- .DW
        001019 => x"0a00", -- .DW
        others => x"0000"  -- NOP
	);
	------------------------------------------------------

begin

	-- Memory Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		MEM_FILE_ACCESS: process(CLK_I)
		begin
			if rising_edge(CLK_I) then
				-- Data Read --
				if (D_EN_I = '1') then -- valid access
					if (word_mode_en_c = true) then -- read data access
						D_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(D_ADR_I(log2_mem_size_c-1 downto 0))));
					else
						D_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(D_ADR_I(log2_mem_size_c downto 1))));
					end if;
				end if;
				-- Instruction Read --
				if (I_EN_I = '1') then
					if (word_mode_en_c = true) then
						I_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(I_ADR_I(log2_mem_size_c-1 downto 0))));
					else
						I_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(I_ADR_I(log2_mem_size_c downto 1))));
					end if;
				end if;
			end if;
		end process MEM_FILE_ACCESS;



end BOOT_MEM_STRUCTURE;
