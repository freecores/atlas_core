-- ########################################################
-- #         << ATLAS Project - Bootloader ROM >>         #
-- # **************************************************** #
-- #  Initialized with boot loader.                       #
-- # **************************************************** #
-- #  Last modified: 14.04.2014                           #
-- # **************************************************** #
-- #  by Stephan Nolting 4788, Hanover, Germany           #
-- ########################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.atlas_core_package.all;

entity BOOT_MEM is
	port	(
				-- Host Interface --
				CLK_I           : in  std_logic; -- global clock line
				I_ADR_I         : in  std_logic_vector(15 downto 0); -- instruction adr
				I_EN_I          : in  std_logic; -- IR update
				I_DAT_O         : out std_logic_vector(15 downto 0); -- instruction out
				D_EN_I          : in  std_logic; -- access enable
				D_RW_I          : in  std_logic; -- read/write
				D_ADR_I         : in  std_logic_vector(15 downto 0); -- data adr
				D_DAT_I         : in  std_logic_vector(15 downto 0); -- data in
				D_DAT_O         : out std_logic_vector(15 downto 0)  -- data out
			);
end BOOT_MEM;

architecture BOOT_MEM_STRUCTURE of BOOT_MEM is

	-- Internal constants(configuration --
	constant mem_size_c      : natural := 2048; -- 2kB
	constant log2_mem_size_c : natural := log2(mem_size_c/2); -- address width (word boundary!)

	-- Memory Type --
	type mem_file_t is array (0 to (mem_size_c/2)-1) of std_logic_vector(15 downto 0); -- word mem!

	-- MEMORY IMAGE (Bootloader Program) --
	------------------------------------------------------
	constant BOOT_MEM_FILE_C : mem_file_t :=
    (
        000000 => x"bc0e", -- B
        000001 => x"bc04", -- B
        000002 => x"bc03", -- B
        000003 => x"bc02", -- B
        000004 => x"bc01", -- B
        000005 => x"c000", -- LDIL
        000006 => x"cc00", -- LDIH
        000007 => x"ec8a", -- MCR
        000008 => x"cc19", -- LDIH
        000009 => x"ed0f", -- MCR
        000010 => x"c528", -- LDIL
        000011 => x"c907", -- LDIH
        000012 => x"be86", -- BL
        000013 => x"bc00", -- B
        000014 => x"ec11", -- MRC
        000015 => x"ec88", -- MCR
        000016 => x"ec8a", -- MCR
        000017 => x"c380", -- LDIL
        000018 => x"cff8", -- LDIH
        000019 => x"1c07", -- STSR
        000020 => x"2800", -- CLR
        000021 => x"ec08", -- MCR
        000022 => x"ec0b", -- MCR
        000023 => x"ec0e", -- MCR
        000024 => x"ec00", -- MRC
        000025 => x"ed88", -- MCR
        000026 => x"c002", -- LDIL
        000027 => x"ed8b", -- MCR
        000028 => x"c064", -- LDIL
        000029 => x"ed8d", -- MCR
        000030 => x"c901", -- LDIH
        000031 => x"ed2f", -- MCR
        000032 => x"ec17", -- MRC
        000033 => x"ec97", -- MRC
        000034 => x"c160", -- LDIL
        000035 => x"c909", -- LDIH
        000036 => x"c18f", -- LDIL
        000037 => x"0923", -- ADD
        000038 => x"29b3", -- CLR
        000039 => x"2a44", -- CLR
        000040 => x"100a", -- SUBS
        000041 => x"149b", -- SBCS
        000042 => x"9003", -- BMI
        000043 => x"0241", -- INC
        000044 => x"bdfc", -- B
        000045 => x"ed49", -- MCR
        000046 => x"ec22", -- MRC
        000047 => x"d406", -- SBR
        000048 => x"ed0a", -- MCR
        000049 => x"c536", -- LDIL
        000050 => x"c905", -- LDIH
        000051 => x"be5f", -- BL
        000052 => x"c12c", -- LDIL
        000053 => x"c906", -- LDIH
        000054 => x"be5c", -- BL
        000055 => x"ee11", -- MRC
        000056 => x"be5e", -- BL
        000057 => x"c13c", -- LDIL
        000058 => x"c906", -- LDIH
        000059 => x"be57", -- BL
        000060 => x"ee97", -- MRC
        000061 => x"ee17", -- MRC
        000062 => x"be58", -- BL
        000063 => x"0250", -- MOV
        000064 => x"be56", -- BL
        000065 => x"be52", -- BL
        000066 => x"ec27", -- MRC
        000067 => x"c083", -- LDIL
        000068 => x"2001", -- AND
        000069 => x"c330", -- LDIL
        000070 => x"0b60", -- ADD
        000071 => x"bc0f", -- B
        000072 => x"c55c", -- LDIL
        000073 => x"c906", -- LDIH
        000074 => x"be48", -- BL
        000075 => x"c14c", -- LDIL
        000076 => x"c907", -- LDIH
        000077 => x"be45", -- BL
        000078 => x"c512", -- LDIL
        000079 => x"c907", -- LDIH
        000080 => x"be42", -- BL
        000081 => x"be44", -- BL
        000082 => x"0300", -- MOV
        000083 => x"0080", -- MOV
        000084 => x"be40", -- BL
        000085 => x"be3e", -- BL
        000086 => x"c0b0", -- LDIL
        000087 => x"181e", -- CMP
        000088 => x"81f0", -- BEQ
        000089 => x"c0b1", -- LDIL
        000090 => x"181e", -- CMP
        000091 => x"809a", -- BEQ
        000092 => x"c0b2", -- LDIL
        000093 => x"181e", -- CMP
        000094 => x"8064", -- BEQ
        000095 => x"c0b3", -- LDIL
        000096 => x"181e", -- CMP
        000097 => x"802b", -- BEQ
        000098 => x"c0b4", -- LDIL
        000099 => x"181e", -- CMP
        000100 => x"8033", -- BEQ
        000101 => x"c0bf", -- LDIL
        000102 => x"181e", -- CMP
        000103 => x"8405", -- BNE
        000104 => x"c102", -- LDIL
        000105 => x"c901", -- LDIH
        000106 => x"be28", -- BL
        000107 => x"bde3", -- B
        000108 => x"c2bc", -- LDIL
        000109 => x"ca83", -- LDIH
        000110 => x"c0f0", -- LDIL
        000111 => x"181e", -- CMP
        000112 => x"f705", -- RBAEQ
        000113 => x"c0e4", -- LDIL
        000114 => x"181e", -- CMP
        000115 => x"80f0", -- BEQ
        000116 => x"c2e2", -- LDIL
        000117 => x"ca85", -- LDIH
        000118 => x"c0f7", -- LDIL
        000119 => x"181e", -- CMP
        000120 => x"f705", -- RBAEQ
        000121 => x"c0f2", -- LDIL
        000122 => x"181e", -- CMP
        000123 => x"85d3", -- BNE
        000124 => x"2800", -- CLR
        000125 => x"c080", -- LDIL
        000126 => x"cc80", -- LDIH
        000127 => x"ec99", -- MCR
        000128 => x"3400", -- GT
        000129 => x"4b65", -- .DW
        000130 => x"6570", -- .DW
        000131 => x"696e", -- .DW
        000132 => x"2720", -- .DW
        000133 => x"6974", -- .DW
        000134 => x"2063", -- .DW
        000135 => x"6f75", -- .DW
        000136 => x"6e74", -- .DW
        000137 => x"7279", -- .DW
        000138 => x"210d", -- .DW
        000139 => x"0a00", -- .DW
        000140 => x"c14c", -- LDIL
        000141 => x"c906", -- LDIH
        000142 => x"be04", -- BL
        000143 => x"2800", -- CLR
        000144 => x"2100", -- STUB
        000145 => x"bca6", -- B
        000146 => x"bc9b", -- B
        000147 => x"bc9b", -- B
        000148 => x"bc9b", -- B
        000149 => x"bc9b", -- B
        000150 => x"bc9e", -- B
        000151 => x"c52c", -- LDIL
        000152 => x"c906", -- LDIH
        000153 => x"be94", -- BL
        000154 => x"be9c", -- BL
        000155 => x"edca", -- MCR
        000156 => x"be9a", -- BL
        000157 => x"edc9", -- MCR
        000158 => x"c424", -- LDIL
        000159 => x"c805", -- LDIH
        000160 => x"3404", -- GTL
        000161 => x"be8d", -- BL
        000162 => x"be93", -- BL
        000163 => x"c47e", -- LDIL
        000164 => x"cc4a", -- LDIH
        000165 => x"180e", -- CMP
        000166 => x"848c", -- BNE
        000167 => x"be8e", -- BL
        000168 => x"3f64", -- SFT
        000169 => x"2066", -- STUB
        000170 => x"be8b", -- BL
        000171 => x"20e6", -- STUB
        000172 => x"be89", -- BL
        000173 => x"2166", -- STUB
        000174 => x"be87", -- BL
        000175 => x"21e6", -- STUB
        000176 => x"be85", -- BL
        000177 => x"2266", -- STUB
        000178 => x"be83", -- BL
        000179 => x"22e6", -- STUB
        000180 => x"be81", -- BL
        000181 => x"2366", -- STUB
        000182 => x"c280", -- LDIL
        000183 => x"ecda", -- MCR
        000184 => x"ec5d", -- MCR
        000185 => x"be7c", -- BL
        000186 => x"7f5a", -- STR
        000187 => x"ec05", -- MRC
        000188 => x"2806", -- EOR
        000189 => x"ec0d", -- MCR
        000190 => x"2400", -- LDUB
        000191 => x"1858", -- CMP
        000192 => x"85f9", -- BNE
        000193 => x"bc59", -- B
        000194 => x"c14c", -- LDIL
        000195 => x"c906", -- LDIH
        000196 => x"be69", -- BL
        000197 => x"c100", -- LDIL
        000198 => x"be28", -- BL
        000199 => x"c47e", -- LDIL
        000200 => x"cc4a", -- LDIH
        000201 => x"180d", -- CMP
        000202 => x"8468", -- BNE
        000203 => x"c102", -- LDIL
        000204 => x"be22", -- BL
        000205 => x"2055", -- STUB
        000206 => x"c104", -- LDIL
        000207 => x"be1f", -- BL
        000208 => x"20d5", -- STUB
        000209 => x"c106", -- LDIL
        000210 => x"be1c", -- BL
        000211 => x"2155", -- STUB
        000212 => x"c108", -- LDIL
        000213 => x"be19", -- BL
        000214 => x"21d5", -- STUB
        000215 => x"c10a", -- LDIL
        000216 => x"be16", -- BL
        000217 => x"2255", -- STUB
        000218 => x"c10c", -- LDIL
        000219 => x"be13", -- BL
        000220 => x"22d5", -- STUB
        000221 => x"c10e", -- LDIL
        000222 => x"be10", -- BL
        000223 => x"2355", -- STUB
        000224 => x"c200", -- LDIL
        000225 => x"ecca", -- MCR
        000226 => x"ec4d", -- MCR
        000227 => x"c010", -- LDIL
        000228 => x"0940", -- ADD
        000229 => x"be09", -- BL
        000230 => x"7eca", -- STR
        000231 => x"ec05", -- MRC
        000232 => x"2805", -- EOR
        000233 => x"ec0d", -- MCR
        000234 => x"2400", -- LDUB
        000235 => x"1848", -- CMP
        000236 => x"85f7", -- BNE
        000237 => x"bc2d", -- B
        000238 => x"0370", -- MOV
        000239 => x"be42", -- BL
        000240 => x"3eb0", -- SFT
        000241 => x"0121", -- INC
        000242 => x"be3f", -- BL
        000243 => x"26d3", -- ORR
        000244 => x"3460", -- RET
        000245 => x"c164", -- LDIL
        000246 => x"c906", -- LDIH
        000247 => x"be36", -- BL
        000248 => x"be38", -- BL
        000249 => x"3c80", -- SFT
        000250 => x"be36", -- BL
        000251 => x"2490", -- ORR
        000252 => x"c47e", -- LDIL
        000253 => x"cc4a", -- LDIH
        000254 => x"1818", -- CMP
        000255 => x"8433", -- BNE
        000256 => x"be27", -- BL
        000257 => x"3c94", -- SFT
        000258 => x"2011", -- STUB
        000259 => x"be24", -- BL
        000260 => x"2091", -- STUB
        000261 => x"be22", -- BL
        000262 => x"2111", -- STUB
        000263 => x"be20", -- BL
        000264 => x"2191", -- STUB
        000265 => x"be1e", -- BL
        000266 => x"2211", -- STUB
        000267 => x"be1c", -- BL
        000268 => x"2291", -- STUB
        000269 => x"be1a", -- BL
        000270 => x"2311", -- STUB
        000271 => x"2ad5", -- CLR
        000272 => x"ecda", -- MCR
        000273 => x"ec5d", -- MCR
        000274 => x"be15", -- BL
        000275 => x"7cda", -- STR
        000276 => x"ec05", -- MRC
        000277 => x"2801", -- EOR
        000278 => x"ec0d", -- MCR
        000279 => x"2400", -- LDUB
        000280 => x"1858", -- CMP
        000281 => x"85f9", -- BNE
        000282 => x"ec11", -- MRC
        000283 => x"ec8a", -- MCR
        000284 => x"c50a", -- LDIL
        000285 => x"c906", -- LDIH
        000286 => x"be0f", -- BL
        000287 => x"ec05", -- MRC
        000288 => x"2491", -- LDUB
        000289 => x"1809", -- CMP
        000290 => x"8015", -- BEQ
        000291 => x"c536", -- LDIL
        000292 => x"c907", -- LDIH
        000293 => x"be08", -- BL
        000294 => x"bccb", -- B
        000295 => x"0370", -- MOV
        000296 => x"be08", -- BL
        000297 => x"3c80", -- SFT
        000298 => x"be06", -- BL
        000299 => x"2490", -- ORR
        000300 => x"3460", -- RET
        000301 => x"bcc7", -- B
        000302 => x"bcd0", -- B
        000303 => x"bcd4", -- B
        000304 => x"bcd8", -- B
        000305 => x"bc6b", -- B
        000306 => x"bcbc", -- B
        000307 => x"bd1b", -- B
        000308 => x"bc69", -- B
        000309 => x"bcbe", -- B
        000310 => x"bcd7", -- B
        000311 => x"c54a", -- LDIL
        000312 => x"c906", -- LDIH
        000313 => x"bebb", -- BL
        000314 => x"ee05", -- MRC
        000315 => x"bef7", -- BL
        000316 => x"bec2", -- BL
        000317 => x"c17a", -- LDIL
        000318 => x"c906", -- LDIH
        000319 => x"beb5", -- BL
        000320 => x"24aa", -- LDUBS
        000321 => x"8010", -- BEQ
        000322 => x"c0a2", -- LDIL
        000323 => x"bec0", -- BL
        000324 => x"24a2", -- LDUB
        000325 => x"be18", -- BL
        000326 => x"24b3", -- LDUB
        000327 => x"be16", -- BL
        000328 => x"24c4", -- LDUB
        000329 => x"be14", -- BL
        000330 => x"24d5", -- LDUB
        000331 => x"be12", -- BL
        000332 => x"24e6", -- LDUB
        000333 => x"be10", -- BL
        000334 => x"c0a2", -- LDIL
        000335 => x"beb4", -- BL
        000336 => x"beae", -- BL
        000337 => x"bead", -- BL
        000338 => x"c080", -- LDIL
        000339 => x"ccc0", -- LDIH
        000340 => x"1c01", -- STSR
        000341 => x"2800", -- CLR
        000342 => x"ed0f", -- MCR
        000343 => x"ec88", -- MCR
        000344 => x"ec8b", -- MCR
        000345 => x"ec8c", -- MCR
        000346 => x"ec8a", -- MCR
        000347 => x"ec89", -- MCR
        000348 => x"3400", -- GT
        000349 => x"0370", -- MOV
        000350 => x"3c90", -- SFT
        000351 => x"bea4", -- BL
        000352 => x"3c90", -- SFT
        000353 => x"bea2", -- BL
        000354 => x"3460", -- RET
        000355 => x"c51e", -- LDIL
        000356 => x"c906", -- LDIH
        000357 => x"be8f", -- BL
        000358 => x"bea7", -- BL
        000359 => x"c524", -- LDIL
        000360 => x"c905", -- LDIH
        000361 => x"3424", -- GTL
        000362 => x"ecca", -- MCR
        000363 => x"be93", -- BL
        000364 => x"c280", -- LDIL
        000365 => x"c00f", -- LDIL
        000366 => x"2058", -- ANDS
        000367 => x"840a", -- BNE
        000368 => x"be8e", -- BL
        000369 => x"c0a4", -- LDIL
        000370 => x"be91", -- BL
        000371 => x"0250", -- MOV
        000372 => x"bebe", -- BL
        000373 => x"c0ba", -- LDIL
        000374 => x"be8d", -- BL
        000375 => x"c0a0", -- LDIL
        000376 => x"be8b", -- BL
        000377 => x"7a5a", -- LDR
        000378 => x"c0a0", -- LDIL
        000379 => x"be88", -- BL
        000380 => x"beb6", -- BL
        000381 => x"c00f", -- LDIL
        000382 => x"2058", -- ANDS
        000383 => x"8414", -- BNE
        000384 => x"c0a0", -- LDIL
        000385 => x"be82", -- BL
        000386 => x"be81", -- BL
        000387 => x"c010", -- LDIL
        000388 => x"1250", -- SUB
        000389 => x"c470", -- LDIL
        000390 => x"2240", -- AND
        000391 => x"78c9", -- LDR
        000392 => x"3c90", -- SFT
        000393 => x"c880", -- LDIH
        000394 => x"c020", -- LDIL
        000395 => x"1818", -- CMP
        000396 => x"a402", -- BLS
        000397 => x"c0ae", -- LDIL
        000398 => x"be75", -- BL
        000399 => x"c08f", -- LDIL
        000400 => x"2014", -- AND
        000401 => x"3409", -- TEQ
        000402 => x"85f5", -- BNE
        000403 => x"ec20", -- MRC
        000404 => x"dc0f", -- STB
        000405 => x"b804", -- BTS
        000406 => x"c5fe", -- LDIL
        000407 => x"343d", -- TEQ
        000408 => x"85d5", -- BNE
        000409 => x"be6f", -- BL
        000410 => x"2800", -- CLR
        000411 => x"3400", -- GT
        000412 => x"bc56", -- B
        000413 => x"bc95", -- B
        000414 => x"c001", -- LDIL
        000415 => x"ed0c", -- MCR
        000416 => x"c050", -- LDIL
        000417 => x"c83f", -- LDIH
        000418 => x"ed0a", -- MCR
        000419 => x"c000", -- LDIL
        000420 => x"c801", -- LDIH
        000421 => x"beab", -- BL
        000422 => x"c156", -- LDIL
        000423 => x"c906", -- LDIH
        000424 => x"be4c", -- BL
        000425 => x"c164", -- LDIL
        000426 => x"c906", -- LDIH
        000427 => x"be49", -- BL
        000428 => x"be5c", -- BL
        000429 => x"3c80", -- SFT
        000430 => x"be5a", -- BL
        000431 => x"2410", -- ORR
        000432 => x"c4fe", -- LDIL
        000433 => x"ccca", -- LDIH
        000434 => x"1809", -- CMP
        000435 => x"843b", -- BNE
        000436 => x"c100", -- LDIL
        000437 => x"c6fe", -- LDIL
        000438 => x"ceca", -- LDIH
        000439 => x"be30", -- BL
        000440 => x"be50", -- BL
        000441 => x"3c80", -- SFT
        000442 => x"be4e", -- BL
        000443 => x"2690", -- ORR
        000444 => x"3ed4", -- SFT
        000445 => x"2055", -- STUB
        000446 => x"c102", -- LDIL
        000447 => x"be28", -- BL
        000448 => x"be48", -- BL
        000449 => x"3c80", -- SFT
        000450 => x"be46", -- BL
        000451 => x"2690", -- ORR
        000452 => x"20d5", -- STUB
        000453 => x"c104", -- LDIL
        000454 => x"be21", -- BL
        000455 => x"c106", -- LDIL
        000456 => x"be40", -- BL
        000457 => x"0180", -- MOV
        000458 => x"be8c", -- BL
        000459 => x"0121", -- INC
        000460 => x"c010", -- LDIL
        000461 => x"1828", -- CMP
        000462 => x"85fa", -- BNE
        000463 => x"c110", -- LDIL
        000464 => x"2ad5", -- CLR
        000465 => x"be37", -- BL
        000466 => x"0180", -- MOV
        000467 => x"be83", -- BL
        000468 => x"0121", -- INC
        000469 => x"2400", -- LDUB
        000470 => x"02d1", -- INC
        000471 => x"1858", -- CMP
        000472 => x"85f9", -- BNE
        000473 => x"c001", -- LDIL
        000474 => x"ed0c", -- MCR
        000475 => x"c050", -- LDIL
        000476 => x"c83f", -- LDIH
        000477 => x"ed0a", -- MCR
        000478 => x"c00c", -- LDIL
        000479 => x"c801", -- LDIH
        000480 => x"be70", -- BL
        000481 => x"c50a", -- LDIL
        000482 => x"c906", -- LDIH
        000483 => x"be11", -- BL
        000484 => x"c690", -- LDIL
        000485 => x"ca80", -- LDIH
        000486 => x"3450", -- GT
        000487 => x"0370", -- MOV
        000488 => x"3dd0", -- SFT
        000489 => x"be6d", -- BL
        000490 => x"0121", -- INC
        000491 => x"01d0", -- MOV
        000492 => x"be6a", -- BL
        000493 => x"3460", -- RET
        000494 => x"c51a", -- LDIL
        000495 => x"c907", -- LDIH
        000496 => x"be04", -- BL
        000497 => x"bcba", -- B
        000498 => x"bc94", -- B
        000499 => x"bca5", -- B
        000500 => x"01f0", -- MOV
        000501 => x"7829", -- LDR
        000502 => x"c080", -- LDIL
        000503 => x"ccff", -- LDIH
        000504 => x"2081", -- AND
        000505 => x"3c98", -- SFTS
        000506 => x"8003", -- BEQ
        000507 => x"be08", -- BL
        000508 => x"bdf9", -- B
        000509 => x"3430", -- RET
        000510 => x"0170", -- MOV
        000511 => x"c08d", -- LDIL
        000512 => x"be03", -- BL
        000513 => x"c08a", -- LDIL
        000514 => x"03a0", -- MOV
        000515 => x"ec22", -- MRC
        000516 => x"dc05", -- STB
        000517 => x"b9fe", -- BTS
        000518 => x"ed18", -- MCR
        000519 => x"3470", -- RET
        000520 => x"ec20", -- MRC
        000521 => x"dc8f", -- STBI
        000522 => x"b9fe", -- BTS
        000523 => x"c800", -- LDIH
        000524 => x"3470", -- RET
        000525 => x"0170", -- MOV
        000526 => x"c200", -- LDIL
        000527 => x"c184", -- LDIL
        000528 => x"bff8", -- BL
        000529 => x"c0c6", -- LDIL
        000530 => x"1809", -- CMP
        000531 => x"9003", -- BMI
        000532 => x"c0a0", -- LDIL
        000533 => x"1001", -- SUB
        000534 => x"c0b0", -- LDIL
        000535 => x"1809", -- CMP
        000536 => x"91f8", -- BMI
        000537 => x"c0c6", -- LDIL
        000538 => x"1818", -- CMP
        000539 => x"91f5", -- BMI
        000540 => x"c0b9", -- LDIL
        000541 => x"1818", -- CMP
        000542 => x"a404", -- BLS
        000543 => x"c0c1", -- LDIL
        000544 => x"1809", -- CMP
        000545 => x"a1ef", -- BHI
        000546 => x"0080", -- MOV
        000547 => x"bfe0", -- BL
        000548 => x"c030", -- LDIL
        000549 => x"1090", -- SUB
        000550 => x"c009", -- LDIL
        000551 => x"1809", -- CMP
        000552 => x"a402", -- BLS
        000553 => x"0497", -- DEC
        000554 => x"3e42", -- SFT
        000555 => x"3e42", -- SFT
        000556 => x"3e42", -- SFT
        000557 => x"3e42", -- SFT
        000558 => x"2641", -- ORR
        000559 => x"05b9", -- DECS
        000560 => x"85e0", -- BNE
        000561 => x"3420", -- RET
        000562 => x"0370", -- MOV
        000563 => x"3d42", -- SFT
        000564 => x"3d22", -- SFT
        000565 => x"3d22", -- SFT
        000566 => x"3d22", -- SFT
        000567 => x"be0f", -- BL
        000568 => x"bfcb", -- BL
        000569 => x"3d40", -- SFT
        000570 => x"be0c", -- BL
        000571 => x"bfc8", -- BL
        000572 => x"3d45", -- SFT
        000573 => x"3d25", -- SFT
        000574 => x"3d25", -- SFT
        000575 => x"3d25", -- SFT
        000576 => x"be06", -- BL
        000577 => x"bfc2", -- BL
        000578 => x"0140", -- MOV
        000579 => x"be03", -- BL
        000580 => x"bfbf", -- BL
        000581 => x"3460", -- RET
        000582 => x"c08f", -- LDIL
        000583 => x"2121", -- AND
        000584 => x"c089", -- LDIL
        000585 => x"181a", -- CMP
        000586 => x"8803", -- BCS
        000587 => x"c0b0", -- LDIL
        000588 => x"bc02", -- B
        000589 => x"c0b7", -- LDIL
        000590 => x"0892", -- ADD
        000591 => x"3470", -- RET
        000592 => x"ed0b", -- MCR
        000593 => x"ec22", -- MRC
        000594 => x"dc03", -- STB
        000595 => x"b9fe", -- BTS
        000596 => x"ec23", -- MRC
        000597 => x"3470", -- RET
        000598 => x"00f0", -- MOV
        000599 => x"c050", -- LDIL
        000600 => x"c837", -- LDIH
        000601 => x"ed0a", -- MCR
        000602 => x"c001", -- LDIL
        000603 => x"ed0c", -- MCR
        000604 => x"c006", -- LDIL
        000605 => x"bff3", -- BL
        000606 => x"c050", -- LDIL
        000607 => x"c83f", -- LDIH
        000608 => x"ed0a", -- MCR
        000609 => x"c000", -- LDIL
        000610 => x"c805", -- LDIH
        000611 => x"bfed", -- BL
        000612 => x"dc01", -- STB
        000613 => x"b805", -- BTS
        000614 => x"c546", -- LDIL
        000615 => x"c907", -- LDIH
        000616 => x"bf8c", -- BL
        000617 => x"bc42", -- B
        000618 => x"c040", -- LDIL
        000619 => x"c83f", -- LDIH
        000620 => x"ed0a", -- MCR
        000621 => x"c001", -- LDIL
        000622 => x"ed0c", -- MCR
        000623 => x"3c20", -- SFT
        000624 => x"c802", -- LDIH
        000625 => x"bfdf", -- BL
        000626 => x"03a0", -- MOV
        000627 => x"cb80", -- LDIH
        000628 => x"3ff0", -- SFT
        000629 => x"0030", -- MOV
        000630 => x"c800", -- LDIH
        000631 => x"2407", -- ORR
        000632 => x"bfd8", -- BL
        000633 => x"2800", -- CLR
        000634 => x"ed0c", -- MCR
        000635 => x"c050", -- LDIL
        000636 => x"c83f", -- LDIH
        000637 => x"ed0a", -- MCR
        000638 => x"c001", -- LDIL
        000639 => x"ed0c", -- MCR
        000640 => x"c000", -- LDIL
        000641 => x"c805", -- LDIH
        000642 => x"bfce", -- BL
        000643 => x"dc00", -- STB
        000644 => x"b9fc", -- BTS
        000645 => x"3410", -- RET
        000646 => x"00f0", -- MOV
        000647 => x"c040", -- LDIL
        000648 => x"c83f", -- LDIH
        000649 => x"ed0a", -- MCR
        000650 => x"c001", -- LDIL
        000651 => x"ed0c", -- MCR
        000652 => x"3c20", -- SFT
        000653 => x"c803", -- LDIH
        000654 => x"bfc2", -- BL
        000655 => x"0020", -- MOV
        000656 => x"c800", -- LDIH
        000657 => x"3c00", -- SFT
        000658 => x"bfbe", -- BL
        000659 => x"29b3", -- CLR
        000660 => x"ed3c", -- MCR
        000661 => x"0180", -- MOV
        000662 => x"c980", -- LDIH
        000663 => x"3410", -- RET
        000664 => x"e5b0", -- CDP
        000665 => x"ec30", -- MRC
        000666 => x"dc06", -- STB
        000667 => x"b9fe", -- BTS
        000668 => x"c306", -- LDIL
        000669 => x"200e", -- ANDS
        000670 => x"840a", -- BNE
        000671 => x"ecb1", -- MRC
        000672 => x"ef32", -- MRC
        000673 => x"2800", -- CLR
        000674 => x"009a", -- INCS
        000675 => x"0f60", -- ADC
        000676 => x"ed99", -- MCR
        000677 => x"edea", -- MCR
        000678 => x"ef34", -- MRC
        000679 => x"3470", -- RET
        000680 => x"c558", -- LDIL
        000681 => x"c907", -- LDIH
        000682 => x"bf4a", -- BL
        000683 => x"c566", -- LDIL
        000684 => x"c907", -- LDIH
        000685 => x"bf47", -- BL
        000686 => x"bf5a", -- BL
        000687 => x"2800", -- CLR
        000688 => x"3400", -- GT
        000689 => x"c52c", -- LDIL
        000690 => x"c906", -- LDIH
        000691 => x"bf41", -- BL
        000692 => x"bf59", -- BL
        000693 => x"edca", -- MCR
        000694 => x"bf57", -- BL
        000695 => x"edc9", -- MCR
        000696 => x"be1a", -- BL
        000697 => x"bf45", -- BL
        000698 => x"c53a", -- LDIL
        000699 => x"c906", -- LDIH
        000700 => x"bf38", -- BL
        000701 => x"bf50", -- BL
        000702 => x"02c0", -- MOV
        000703 => x"be13", -- BL
        000704 => x"345d", -- TEQ
        000705 => x"800d", -- BEQ
        000706 => x"06d1", -- DEC
        000707 => x"bf3b", -- BL
        000708 => x"bfd4", -- BL
        000709 => x"c556", -- LDIL
        000710 => x"c906", -- LDIH
        000711 => x"bf2d", -- BL
        000712 => x"0260", -- MOV
        000713 => x"bf69", -- BL
        000714 => x"eca0", -- MRC
        000715 => x"dc1f", -- STB
        000716 => x"b802", -- BTS
        000717 => x"bdf3", -- B
        000718 => x"bf30", -- BL
        000719 => x"c69c", -- LDIL
        000720 => x"ca80", -- LDIH
        000721 => x"3450", -- GT
        000722 => x"0170", -- MOV
        000723 => x"bf35", -- BL
        000724 => x"c08d", -- LDIL
        000725 => x"1809", -- CMP
        000726 => x"f702", -- RBAEQ
        000727 => x"c088", -- LDIL
        000728 => x"1809", -- CMP
        000729 => x"81f5", -- BEQ
        000730 => x"bdf9", -- B
        000731 => x"0d0a", -- .DW
        000732 => x"0d0a", -- .DW
        000733 => x"4174", -- .DW
        000734 => x"6c61", -- .DW
        000735 => x"732d", -- .DW
        000736 => x"324b", -- .DW
        000737 => x"2042", -- .DW
        000738 => x"6f6f", -- .DW
        000739 => x"746c", -- .DW
        000740 => x"6f61", -- .DW
        000741 => x"6465", -- .DW
        000742 => x"7220", -- .DW
        000743 => x"2d20", -- .DW
        000744 => x"5632", -- .DW
        000745 => x"3031", -- .DW
        000746 => x"3430", -- .DW
        000747 => x"3431", -- .DW
        000748 => x"340d", -- .DW
        000749 => x"0a62", -- .DW
        000750 => x"7920", -- .DW
        000751 => x"5374", -- .DW
        000752 => x"6570", -- .DW
        000753 => x"6861", -- .DW
        000754 => x"6e20", -- .DW
        000755 => x"4e6f", -- .DW
        000756 => x"6c74", -- .DW
        000757 => x"696e", -- .DW
        000758 => x"672c", -- .DW
        000759 => x"2073", -- .DW
        000760 => x"746e", -- .DW
        000761 => x"6f6c", -- .DW
        000762 => x"7469", -- .DW
        000763 => x"6e67", -- .DW
        000764 => x"4067", -- .DW
        000765 => x"6d61", -- .DW
        000766 => x"696c", -- .DW
        000767 => x"2e63", -- .DW
        000768 => x"6f6d", -- .DW
        000769 => x"0d0a", -- .DW
        000770 => x"7777", -- .DW
        000771 => x"772e", -- .DW
        000772 => x"6f70", -- .DW
        000773 => x"656e", -- .DW
        000774 => x"636f", -- .DW
        000775 => x"7265", -- .DW
        000776 => x"732e", -- .DW
        000777 => x"6f72", -- .DW
        000778 => x"672f", -- .DW
        000779 => x"7072", -- .DW
        000780 => x"6f6a", -- .DW
        000781 => x"6563", -- .DW
        000782 => x"742c", -- .DW
        000783 => x"6174", -- .DW
        000784 => x"6c61", -- .DW
        000785 => x"735f", -- .DW
        000786 => x"636f", -- .DW
        000787 => x"7265", -- .DW
        000788 => x"0d0a", -- .DW
        000789 => x"0000", -- .DW
        000790 => x"0d0a", -- .DW
        000791 => x"426f", -- .DW
        000792 => x"6f74", -- .DW
        000793 => x"2070", -- .DW
        000794 => x"6167", -- .DW
        000795 => x"653a", -- .DW
        000796 => x"2030", -- .DW
        000797 => x"7800", -- .DW
        000798 => x"0d0a", -- .DW
        000799 => x"436c", -- .DW
        000800 => x"6f63", -- .DW
        000801 => x"6b28", -- .DW
        000802 => x"487a", -- .DW
        000803 => x"293a", -- .DW
        000804 => x"2030", -- .DW
        000805 => x"7800", -- .DW
        000806 => x"426f", -- .DW
        000807 => x"6f74", -- .DW
        000808 => x"696e", -- .DW
        000809 => x"670d", -- .DW
        000810 => x"0a00", -- .DW
        000811 => x"4275", -- .DW
        000812 => x"726e", -- .DW
        000813 => x"2045", -- .DW
        000814 => x"4550", -- .DW
        000815 => x"524f", -- .DW
        000816 => x"4d0d", -- .DW
        000817 => x"0a00", -- .DW
        000818 => x"5761", -- .DW
        000819 => x"6974", -- .DW
        000820 => x"696e", -- .DW
        000821 => x"6720", -- .DW
        000822 => x"666f", -- .DW
        000823 => x"7220", -- .DW
        000824 => x"6461", -- .DW
        000825 => x"7461", -- .DW
        000826 => x"2e2e", -- .DW
        000827 => x"2e0d", -- .DW
        000828 => x"0a00", -- .DW
        000829 => x"5374", -- .DW
        000830 => x"6172", -- .DW
        000831 => x"7469", -- .DW
        000832 => x"6e67", -- .DW
        000833 => x"2069", -- .DW
        000834 => x"6d61", -- .DW
        000835 => x"6765", -- .DW
        000836 => x"2000", -- .DW
        000837 => x"446f", -- .DW
        000838 => x"776e", -- .DW
        000839 => x"6c6f", -- .DW
        000840 => x"6164", -- .DW
        000841 => x"2063", -- .DW
        000842 => x"6f6d", -- .DW
        000843 => x"706c", -- .DW
        000844 => x"6574", -- .DW
        000845 => x"650d", -- .DW
        000846 => x"0a00", -- .DW
        000847 => x"5061", -- .DW
        000848 => x"6765", -- .DW
        000849 => x"2028", -- .DW
        000850 => x"3468", -- .DW
        000851 => x"293a", -- .DW
        000852 => x"2024", -- .DW
        000853 => x"0000", -- .DW
        000854 => x"4164", -- .DW
        000855 => x"6472", -- .DW
        000856 => x"2028", -- .DW
        000857 => x"3868", -- .DW
        000858 => x"293a", -- .DW
        000859 => x"2024", -- .DW
        000860 => x"0000", -- .DW
        000861 => x"2377", -- .DW
        000862 => x"6f72", -- .DW
        000863 => x"6473", -- .DW
        000864 => x"2028", -- .DW
        000865 => x"3468", -- .DW
        000866 => x"293a", -- .DW
        000867 => x"2024", -- .DW
        000868 => x"0000", -- .DW
        000869 => x"4368", -- .DW
        000870 => x"6563", -- .DW
        000871 => x"6b73", -- .DW
        000872 => x"756d", -- .DW
        000873 => x"3a20", -- .DW
        000874 => x"2400", -- .DW
        000875 => x"202d", -- .DW
        000876 => x"3e20", -- .DW
        000877 => x"2400", -- .DW
        000878 => x"0d0a", -- .DW
        000879 => x"636d", -- .DW
        000880 => x"642f", -- .DW
        000881 => x"626f", -- .DW
        000882 => x"6f74", -- .DW
        000883 => x"2d73", -- .DW
        000884 => x"7769", -- .DW
        000885 => x"7463", -- .DW
        000886 => x"683a", -- .DW
        000887 => x"0d0a", -- .DW
        000888 => x"2030", -- .DW
        000889 => x"2f27", -- .DW
        000890 => x"3030", -- .DW
        000891 => x"273a", -- .DW
        000892 => x"2052", -- .DW
        000893 => x"6573", -- .DW
        000894 => x"7461", -- .DW
        000895 => x"7274", -- .DW
        000896 => x"2063", -- .DW
        000897 => x"6f6e", -- .DW
        000898 => x"736f", -- .DW
        000899 => x"6c65", -- .DW
        000900 => x"0d0a", -- .DW
        000901 => x"2031", -- .DW
        000902 => x"2f27", -- .DW
        000903 => x"3031", -- .DW
        000904 => x"273a", -- .DW
        000905 => x"2042", -- .DW
        000906 => x"6f6f", -- .DW
        000907 => x"7420", -- .DW
        000908 => x"5541", -- .DW
        000909 => x"5254", -- .DW
        000910 => x"0d0a", -- .DW
        000911 => x"2032", -- .DW
        000912 => x"2f27", -- .DW
        000913 => x"3130", -- .DW
        000914 => x"273a", -- .DW
        000915 => x"2042", -- .DW
        000916 => x"6f6f", -- .DW
        000917 => x"7420", -- .DW
        000918 => x"4545", -- .DW
        000919 => x"5052", -- .DW
        000920 => x"4f4d", -- .DW
        000921 => x"0d0a", -- .DW
        000922 => x"2033", -- .DW
        000923 => x"2f27", -- .DW
        000924 => x"3131", -- .DW
        000925 => x"273a", -- .DW
        000926 => x"2042", -- .DW
        000927 => x"6f6f", -- .DW
        000928 => x"7420", -- .DW
        000929 => x"6d65", -- .DW
        000930 => x"6d6f", -- .DW
        000931 => x"7279", -- .DW
        000932 => x"0d0a", -- .DW
        000933 => x"0000", -- .DW
        000934 => x"2034", -- .DW
        000935 => x"3a20", -- .DW
        000936 => x"426f", -- .DW
        000937 => x"6f74", -- .DW
        000938 => x"2057", -- .DW
        000939 => x"420d", -- .DW
        000940 => x"0a20", -- .DW
        000941 => x"703a", -- .DW
        000942 => x"2042", -- .DW
        000943 => x"7572", -- .DW
        000944 => x"6e20", -- .DW
        000945 => x"4545", -- .DW
        000946 => x"5052", -- .DW
        000947 => x"4f4d", -- .DW
        000948 => x"0d0a", -- .DW
        000949 => x"2064", -- .DW
        000950 => x"3a20", -- .DW
        000951 => x"5241", -- .DW
        000952 => x"4d20", -- .DW
        000953 => x"6475", -- .DW
        000954 => x"6d70", -- .DW
        000955 => x"0d0a", -- .DW
        000956 => x"2072", -- .DW
        000957 => x"3a20", -- .DW
        000958 => x"5265", -- .DW
        000959 => x"7365", -- .DW
        000960 => x"740d", -- .DW
        000961 => x"0a20", -- .DW
        000962 => x"773a", -- .DW
        000963 => x"2057", -- .DW
        000964 => x"4220", -- .DW
        000965 => x"6475", -- .DW
        000966 => x"6d70", -- .DW
        000967 => x"0d0a", -- .DW
        000968 => x"0000", -- .DW
        000969 => x"636d", -- .DW
        000970 => x"643a", -- .DW
        000971 => x"3e20", -- .DW
        000972 => x"0000", -- .DW
        000973 => x"494d", -- .DW
        000974 => x"4147", -- .DW
        000975 => x"4520", -- .DW
        000976 => x"4552", -- .DW
        000977 => x"5221", -- .DW
        000978 => x"0d0a", -- .DW
        000979 => x"0000", -- .DW
        000980 => x"0d0a", -- .DW
        000981 => x"4952", -- .DW
        000982 => x"5120", -- .DW
        000983 => x"4552", -- .DW
        000984 => x"5221", -- .DW
        000985 => x"0d0a", -- .DW
        000986 => x"0000", -- .DW
        000987 => x"4348", -- .DW
        000988 => x"4543", -- .DW
        000989 => x"4b53", -- .DW
        000990 => x"554d", -- .DW
        000991 => x"2045", -- .DW
        000992 => x"5252", -- .DW
        000993 => x"210d", -- .DW
        000994 => x"0a00", -- .DW
        000995 => x"5350", -- .DW
        000996 => x"492f", -- .DW
        000997 => x"4545", -- .DW
        000998 => x"5052", -- .DW
        000999 => x"4f4d", -- .DW
        001000 => x"2045", -- .DW
        001001 => x"5252", -- .DW
        001002 => x"210d", -- .DW
        001003 => x"0a00", -- .DW
        001004 => x"5742", -- .DW
        001005 => x"2042", -- .DW
        001006 => x"5553", -- .DW
        001007 => x"2045", -- .DW
        001008 => x"5252", -- .DW
        001009 => x"210d", -- .DW
        001010 => x"0a00", -- .DW
        001011 => x"5072", -- .DW
        001012 => x"6573", -- .DW
        001013 => x"7320", -- .DW
        001014 => x"616e", -- .DW
        001015 => x"7920", -- .DW
        001016 => x"6b65", -- .DW
        001017 => x"790d", -- .DW
        001018 => x"0a00", -- .DW
        others => x"0000"  -- NOP
	);
	------------------------------------------------------

begin

	-- Memory Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		MEM_FILE_ACCESS: process(CLK_I)
		begin
			if rising_edge(CLK_I) then
				-- Data Read --
				if (D_EN_I = '1') then -- valid access
					if (word_mode_en_c = true) then -- read data access
						D_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(D_ADR_I(log2_mem_size_c-1 downto 0))));
					else
						D_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(D_ADR_I(log2_mem_size_c downto 1))));
					end if;
				end if;
				-- Instruction Read --
				if (I_EN_I = '1') then
					if (word_mode_en_c = true) then
						I_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(I_ADR_I(log2_mem_size_c-1 downto 0))));
					else
						I_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(I_ADR_I(log2_mem_size_c downto 1))));
					end if;
				end if;
			end if;
		end process MEM_FILE_ACCESS;



end BOOT_MEM_STRUCTURE;
