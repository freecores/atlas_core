-- ########################################################
-- #         << ATLAS Project - Bootloader ROM >>         #
-- # **************************************************** #
-- #  Initialized with boot loader.                       #
-- # **************************************************** #
-- #  Last modified: 10.04.2014                           #
-- # **************************************************** #
-- #  by Stephan Nolting 4788, Hanover, Germany           #
-- ########################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.atlas_core_package.all;

entity BOOT_MEM is
	port	(
				-- Host Interface --
				CLK_I           : in  std_logic; -- global clock line
				I_ADR_I         : in  std_logic_vector(15 downto 0); -- instruction adr
				I_EN_I          : in  std_logic; -- IR update
				I_DAT_O         : out std_logic_vector(15 downto 0); -- instruction out
				D_EN_I          : in  std_logic; -- access enable
				D_RW_I          : in  std_logic; -- read/write
				D_ADR_I         : in  std_logic_vector(15 downto 0); -- data adr
				D_DAT_I         : in  std_logic_vector(15 downto 0); -- data in
				D_DAT_O         : out std_logic_vector(15 downto 0)  -- data out
			);
end BOOT_MEM;

architecture BOOT_MEM_STRUCTURE of BOOT_MEM is

	-- Internal constants(configuration --
	constant mem_size_c      : natural := 2048; -- 2kB
	constant log2_mem_size_c : natural := log2(mem_size_c/2); -- address width (word boundary!)

	-- Memory Type --
	type mem_file_t is array (0 to (mem_size_c/2)-1) of std_logic_vector(15 downto 0); -- word mem!

	-- MEMORY IMAGE (Bootloader Program) --
	------------------------------------------------------
	constant BOOT_MEM_FILE_C : mem_file_t :=
    (
    000000 => x"bc0e", -- B
    000001 => x"bc04", -- B
    000002 => x"bc03", -- B
    000003 => x"bc02", -- B
    000004 => x"bc01", -- B
    000005 => x"c000", -- LDIL
    000006 => x"cc00", -- LDIH
    000007 => x"ec8a", -- MCR
    000008 => x"cc19", -- LDIH
    000009 => x"ed0f", -- MCR
    000010 => x"c53a", -- LDIL
    000011 => x"c907", -- LDIH
    000012 => x"be85", -- BL
    000013 => x"bc00", -- B
    000014 => x"ec11", -- MRC
    000015 => x"ec88", -- MCR
    000016 => x"ec8a", -- MCR
    000017 => x"c000", -- LDIL
    000018 => x"ec0b", -- MCR
    000019 => x"ec0e", -- MCR
    000020 => x"c802", -- LDIH
    000021 => x"ec08", -- MCR
    000022 => x"c47f", -- LDIL
    000023 => x"ec09", -- MCR
    000024 => x"ec00", -- MRC
    000025 => x"c080", -- LDIL
    000026 => x"ccf8", -- LDIH
    000027 => x"1c01", -- STSR
    000028 => x"c030", -- LDIL
    000029 => x"c800", -- LDIH
    000030 => x"ed88", -- MCR
    000031 => x"c002", -- LDIL
    000032 => x"ed8b", -- MCR
    000033 => x"c064", -- LDIL
    000034 => x"ed8d", -- MCR
    000035 => x"c801", -- LDIH
    000036 => x"ed0f", -- MCR
    000037 => x"ec17", -- MRC
    000038 => x"ec97", -- MRC
    000039 => x"c160", -- LDIL
    000040 => x"c909", -- LDIH
    000041 => x"c18f", -- LDIL
    000042 => x"0923", -- ADD
    000043 => x"29b3", -- CLR
    000044 => x"2a44", -- CLR
    000045 => x"100a", -- SUBS
    000046 => x"149b", -- SBCS
    000047 => x"9003", -- BMI
    000048 => x"0241", -- INC
    000049 => x"bdfc", -- B
    000050 => x"ed49", -- MCR
    000051 => x"ec22", -- MRC
    000052 => x"d406", -- SBR
    000053 => x"ed0a", -- MCR
    000054 => x"be5d", -- BL
    000055 => x"be5c", -- BL
    000056 => x"c54c", -- LDIL
    000057 => x"c905", -- LDIH
    000058 => x"be57", -- BL
    000059 => x"c13e", -- LDIL
    000060 => x"c906", -- LDIH
    000061 => x"be55", -- BL
    000062 => x"ee11", -- MRC
    000063 => x"be57", -- BL
    000064 => x"be53", -- BL
    000065 => x"c14e", -- LDIL
    000066 => x"c906", -- LDIH
    000067 => x"be4f", -- BL
    000068 => x"ee97", -- MRC
    000069 => x"ee17", -- MRC
    000070 => x"be50", -- BL
    000071 => x"0250", -- MOV
    000072 => x"be4e", -- BL
    000073 => x"be4a", -- BL
    000074 => x"ec27", -- MRC
    000075 => x"c083", -- LDIL
    000076 => x"2001", -- AND
    000077 => x"c330", -- LDIL
    000078 => x"0b60", -- ADD
    000079 => x"bc1c", -- B
    000080 => x"be43", -- BL
    000081 => x"c57a", -- LDIL
    000082 => x"c906", -- LDIH
    000083 => x"be3e", -- BL
    000084 => x"c10a", -- LDIL
    000085 => x"c907", -- LDIH
    000086 => x"be3b", -- BL
    000087 => x"c172", -- LDIL
    000088 => x"c907", -- LDIH
    000089 => x"be38", -- BL
    000090 => x"c502", -- LDIL
    000091 => x"c907", -- LDIH
    000092 => x"be35", -- BL
    000093 => x"c510", -- LDIL
    000094 => x"c907", -- LDIH
    000095 => x"be32", -- BL
    000096 => x"c51a", -- LDIL
    000097 => x"c907", -- LDIH
    000098 => x"be2f", -- BL
    000099 => x"c526", -- LDIL
    000100 => x"c907", -- LDIH
    000101 => x"be2d", -- BL
    000102 => x"be2f", -- BL
    000103 => x"0300", -- MOV
    000104 => x"00e0", -- MOV
    000105 => x"be2b", -- BL
    000106 => x"be29", -- BL
    000107 => x"c0b0", -- LDIL
    000108 => x"181e", -- CMP
    000109 => x"81e3", -- BEQ
    000110 => x"c0b1", -- LDIL
    000111 => x"181e", -- CMP
    000112 => x"8078", -- BEQ
    000113 => x"c0b2", -- LDIL
    000114 => x"181e", -- CMP
    000115 => x"8024", -- BEQ
    000116 => x"c0b3", -- LDIL
    000117 => x"181e", -- CMP
    000118 => x"8015", -- BEQ
    000119 => x"c2f4", -- LDIL
    000120 => x"ca83", -- LDIH
    000121 => x"c0f0", -- LDIL
    000122 => x"181e", -- CMP
    000123 => x"f705", -- RBAEQ
    000124 => x"c6f2", -- LDIL
    000125 => x"ca82", -- LDIH
    000126 => x"c0e4", -- LDIL
    000127 => x"181e", -- CMP
    000128 => x"f705", -- RBAEQ
    000129 => x"c68c", -- LDIL
    000130 => x"ca85", -- LDIH
    000131 => x"c0f7", -- LDIL
    000132 => x"181e", -- CMP
    000133 => x"f705", -- RBAEQ
    000134 => x"c0f2", -- LDIL
    000135 => x"181e", -- CMP
    000136 => x"85db", -- BNE
    000137 => x"2800", -- CLR
    000138 => x"3400", -- GT
    000139 => x"c15e", -- LDIL
    000140 => x"c906", -- LDIH
    000141 => x"be04", -- BL
    000142 => x"2800", -- CLR
    000143 => x"2100", -- STUB
    000144 => x"bcb3", -- B
    000145 => x"bca9", -- B
    000146 => x"bca9", -- B
    000147 => x"bca9", -- B
    000148 => x"bca9", -- B
    000149 => x"bca9", -- B
    000150 => x"bcac", -- B
    000151 => x"c15e", -- LDIL
    000152 => x"c906", -- LDIH
    000153 => x"bea1", -- BL
    000154 => x"c100", -- LDIL
    000155 => x"bea4", -- BL
    000156 => x"3eb0", -- SFT
    000157 => x"c101", -- LDIL
    000158 => x"bea1", -- BL
    000159 => x"26d3", -- ORR
    000160 => x"c47e", -- LDIL
    000161 => x"cc4a", -- LDIH
    000162 => x"180d", -- CMP
    000163 => x"849d", -- BNE
    000164 => x"c102", -- LDIL
    000165 => x"be9a", -- BL
    000166 => x"3eb0", -- SFT
    000167 => x"c103", -- LDIL
    000168 => x"be97", -- BL
    000169 => x"26d3", -- ORR
    000170 => x"2055", -- STUB
    000171 => x"c104", -- LDIL
    000172 => x"be93", -- BL
    000173 => x"3eb0", -- SFT
    000174 => x"c105", -- LDIL
    000175 => x"be90", -- BL
    000176 => x"26d3", -- ORR
    000177 => x"20d5", -- STUB
    000178 => x"c106", -- LDIL
    000179 => x"be8c", -- BL
    000180 => x"3eb0", -- SFT
    000181 => x"c107", -- LDIL
    000182 => x"be89", -- BL
    000183 => x"26d3", -- ORR
    000184 => x"2155", -- STUB
    000185 => x"c108", -- LDIL
    000186 => x"be85", -- BL
    000187 => x"3eb0", -- SFT
    000188 => x"c109", -- LDIL
    000189 => x"be82", -- BL
    000190 => x"26d3", -- ORR
    000191 => x"21d5", -- STUB
    000192 => x"c10a", -- LDIL
    000193 => x"be7e", -- BL
    000194 => x"3eb0", -- SFT
    000195 => x"c10b", -- LDIL
    000196 => x"be7b", -- BL
    000197 => x"26d3", -- ORR
    000198 => x"2255", -- STUB
    000199 => x"c10c", -- LDIL
    000200 => x"be77", -- BL
    000201 => x"3eb0", -- SFT
    000202 => x"c10d", -- LDIL
    000203 => x"be74", -- BL
    000204 => x"26d3", -- ORR
    000205 => x"22d5", -- STUB
    000206 => x"c10e", -- LDIL
    000207 => x"be70", -- BL
    000208 => x"3eb0", -- SFT
    000209 => x"c10f", -- LDIL
    000210 => x"be6d", -- BL
    000211 => x"26d3", -- ORR
    000212 => x"2355", -- STUB
    000213 => x"c300", -- LDIL
    000214 => x"ecea", -- MCR
    000215 => x"23e6", -- STUB
    000216 => x"c010", -- LDIL
    000217 => x"0960", -- ADD
    000218 => x"be65", -- BL
    000219 => x"3eb0", -- SFT
    000220 => x"c011", -- LDIL
    000221 => x"0960", -- ADD
    000222 => x"be61", -- BL
    000223 => x"26d3", -- ORR
    000224 => x"7eea", -- STR
    000225 => x"2477", -- LDUB
    000226 => x"2805", -- EOR
    000227 => x"2380", -- STUB
    000228 => x"2400", -- LDUB
    000229 => x"1868", -- CMP
    000230 => x"85f2", -- BNE
    000231 => x"bc41", -- B
    000232 => x"c15e", -- LDIL
    000233 => x"c906", -- LDIH
    000234 => x"be50", -- BL
    000235 => x"c17a", -- LDIL
    000236 => x"c906", -- LDIH
    000237 => x"be4d", -- BL
    000238 => x"be50", -- BL
    000239 => x"3c80", -- SFT
    000240 => x"be4e", -- BL
    000241 => x"2490", -- ORR
    000242 => x"c47e", -- LDIL
    000243 => x"cc4a", -- LDIH
    000244 => x"1818", -- CMP
    000245 => x"844b", -- BNE
    000246 => x"be48", -- BL
    000247 => x"3c80", -- SFT
    000248 => x"be46", -- BL
    000249 => x"2490", -- ORR
    000250 => x"3c94", -- SFT
    000251 => x"2011", -- STUB
    000252 => x"be42", -- BL
    000253 => x"3c80", -- SFT
    000254 => x"be40", -- BL
    000255 => x"2490", -- ORR
    000256 => x"2091", -- STUB
    000257 => x"be3d", -- BL
    000258 => x"3c80", -- SFT
    000259 => x"be3b", -- BL
    000260 => x"2490", -- ORR
    000261 => x"2111", -- STUB
    000262 => x"be38", -- BL
    000263 => x"3c80", -- SFT
    000264 => x"be36", -- BL
    000265 => x"2490", -- ORR
    000266 => x"2191", -- STUB
    000267 => x"be33", -- BL
    000268 => x"3c80", -- SFT
    000269 => x"be31", -- BL
    000270 => x"2490", -- ORR
    000271 => x"2211", -- STUB
    000272 => x"be2e", -- BL
    000273 => x"3c80", -- SFT
    000274 => x"be2c", -- BL
    000275 => x"2490", -- ORR
    000276 => x"2291", -- STUB
    000277 => x"be29", -- BL
    000278 => x"3c80", -- SFT
    000279 => x"be27", -- BL
    000280 => x"2490", -- ORR
    000281 => x"2311", -- STUB
    000282 => x"2ad5", -- CLR
    000283 => x"ecda", -- MCR
    000284 => x"23d5", -- STUB
    000285 => x"be21", -- BL
    000286 => x"3c80", -- SFT
    000287 => x"be1f", -- BL
    000288 => x"2490", -- ORR
    000289 => x"7cda", -- STR
    000290 => x"2477", -- LDUB
    000291 => x"2801", -- EOR
    000292 => x"2380", -- STUB
    000293 => x"2400", -- LDUB
    000294 => x"1858", -- CMP
    000295 => x"85f6", -- BNE
    000296 => x"ec11", -- MRC
    000297 => x"ec8a", -- MCR
    000298 => x"c524", -- LDIL
    000299 => x"c906", -- LDIH
    000300 => x"be0e", -- BL
    000301 => x"2477", -- LDUB
    000302 => x"2491", -- LDUB
    000303 => x"1809", -- CMP
    000304 => x"8013", -- BEQ
    000305 => x"c546", -- LDIL
    000306 => x"c907", -- LDIH
    000307 => x"be07", -- BL
    000308 => x"c564", -- LDIL
    000309 => x"c907", -- LDIH
    000310 => x"be04", -- BL
    000311 => x"be07", -- BL
    000312 => x"2800", -- CLR
    000313 => x"3400", -- GT
    000314 => x"bcdd", -- B
    000315 => x"bcdf", -- B
    000316 => x"bceb", -- B
    000317 => x"bcef", -- B
    000318 => x"bcf3", -- B
    000319 => x"bc79", -- B
    000320 => x"bccd", -- B
    000321 => x"bd22", -- B
    000322 => x"bc77", -- B
    000323 => x"c514", -- LDIL
    000324 => x"c906", -- LDIH
    000325 => x"bed5", -- BL
    000326 => x"24aa", -- LDUBS
    000327 => x"8024", -- BEQ
    000328 => x"c0a2", -- LDIL
    000329 => x"bee3", -- BL
    000330 => x"24a2", -- LDUB
    000331 => x"3c90", -- SFT
    000332 => x"bee0", -- BL
    000333 => x"3c90", -- SFT
    000334 => x"bede", -- BL
    000335 => x"24b3", -- LDUB
    000336 => x"3c90", -- SFT
    000337 => x"bedb", -- BL
    000338 => x"3c90", -- SFT
    000339 => x"bed9", -- BL
    000340 => x"24c4", -- LDUB
    000341 => x"3c90", -- SFT
    000342 => x"bed6", -- BL
    000343 => x"3c90", -- SFT
    000344 => x"bed4", -- BL
    000345 => x"24d5", -- LDUB
    000346 => x"3c90", -- SFT
    000347 => x"bed1", -- BL
    000348 => x"3c90", -- SFT
    000349 => x"becf", -- BL
    000350 => x"24e6", -- LDUB
    000351 => x"3c90", -- SFT
    000352 => x"becc", -- BL
    000353 => x"3c90", -- SFT
    000354 => x"beca", -- BL
    000355 => x"c0a2", -- LDIL
    000356 => x"bec8", -- BL
    000357 => x"bec2", -- BL
    000358 => x"c564", -- LDIL
    000359 => x"c906", -- LDIH
    000360 => x"beb2", -- BL
    000361 => x"2677", -- LDUB
    000362 => x"be4f", -- BL
    000363 => x"bebc", -- BL
    000364 => x"bebb", -- BL
    000365 => x"2800", -- CLR
    000366 => x"d58e", -- SBR
    000367 => x"d5bf", -- SBR
    000368 => x"1c03", -- STSR
    000369 => x"ed0f", -- MCR
    000370 => x"ec88", -- MCR
    000371 => x"ec88", -- MCR
    000372 => x"ec8b", -- MCR
    000373 => x"ec8c", -- MCR
    000374 => x"ec8a", -- MCR
    000375 => x"ec89", -- MCR
    000376 => x"3400", -- GT
    000377 => x"c538", -- LDIL
    000378 => x"c906", -- LDIH
    000379 => x"be9f", -- BL
    000380 => x"beba", -- BL
    000381 => x"beb4", -- BL
    000382 => x"c08d", -- LDIL
    000383 => x"1809", -- CMP
    000384 => x"8006", -- BEQ
    000385 => x"c088", -- LDIL
    000386 => x"1809", -- CMP
    000387 => x"85fa", -- BNE
    000388 => x"bea3", -- BL
    000389 => x"bdbc", -- B
    000390 => x"ecca", -- MCR
    000391 => x"bea0", -- BL
    000392 => x"c280", -- LDIL
    000393 => x"c00f", -- LDIL
    000394 => x"2058", -- ANDS
    000395 => x"840a", -- BNE
    000396 => x"be9b", -- BL
    000397 => x"c0a4", -- LDIL
    000398 => x"be9e", -- BL
    000399 => x"0250", -- MOV
    000400 => x"becb", -- BL
    000401 => x"c0ba", -- LDIL
    000402 => x"be9a", -- BL
    000403 => x"c0a0", -- LDIL
    000404 => x"be98", -- BL
    000405 => x"7a5a", -- LDR
    000406 => x"c0a0", -- LDIL
    000407 => x"be95", -- BL
    000408 => x"bec3", -- BL
    000409 => x"c00f", -- LDIL
    000410 => x"2058", -- ANDS
    000411 => x"8414", -- BNE
    000412 => x"c0a0", -- LDIL
    000413 => x"be8f", -- BL
    000414 => x"be8e", -- BL
    000415 => x"c010", -- LDIL
    000416 => x"1250", -- SUB
    000417 => x"c470", -- LDIL
    000418 => x"2240", -- AND
    000419 => x"78c9", -- LDR
    000420 => x"3c90", -- SFT
    000421 => x"c880", -- LDIH
    000422 => x"c020", -- LDIL
    000423 => x"1818", -- CMP
    000424 => x"a402", -- BLS
    000425 => x"c0ae", -- LDIL
    000426 => x"be82", -- BL
    000427 => x"c08f", -- LDIL
    000428 => x"2014", -- AND
    000429 => x"3409", -- TEQ
    000430 => x"85f5", -- BNE
    000431 => x"ec20", -- MRC
    000432 => x"dc0f", -- STB
    000433 => x"b804", -- BTS
    000434 => x"c5fe", -- LDIL
    000435 => x"343d", -- TEQ
    000436 => x"85d5", -- BNE
    000437 => x"be7c", -- BL
    000438 => x"2800", -- CLR
    000439 => x"3400", -- GT
    000440 => x"bc5e", -- B
    000441 => x"bca2", -- B
    000442 => x"c001", -- LDIL
    000443 => x"ed0c", -- MCR
    000444 => x"c050", -- LDIL
    000445 => x"c83f", -- LDIH
    000446 => x"ed0a", -- MCR
    000447 => x"c000", -- LDIL
    000448 => x"c801", -- LDIH
    000449 => x"beb8", -- BL
    000450 => x"c16a", -- LDIL
    000451 => x"c906", -- LDIH
    000452 => x"be53", -- BL
    000453 => x"c17a", -- LDIL
    000454 => x"c906", -- LDIH
    000455 => x"be50", -- BL
    000456 => x"be69", -- BL
    000457 => x"3c80", -- SFT
    000458 => x"be67", -- BL
    000459 => x"2410", -- ORR
    000460 => x"c4fe", -- LDIL
    000461 => x"ccca", -- LDIH
    000462 => x"1809", -- CMP
    000463 => x"843e", -- BNE
    000464 => x"c100", -- LDIL
    000465 => x"c5ca", -- LDIL
    000466 => x"bead", -- BL
    000467 => x"c101", -- LDIL
    000468 => x"c5fe", -- LDIL
    000469 => x"beaa", -- BL
    000470 => x"be5b", -- BL
    000471 => x"3c80", -- SFT
    000472 => x"be59", -- BL
    000473 => x"2690", -- ORR
    000474 => x"3ed4", -- SFT
    000475 => x"2055", -- STUB
    000476 => x"c102", -- LDIL
    000477 => x"3dd0", -- SFT
    000478 => x"bea1", -- BL
    000479 => x"c103", -- LDIL
    000480 => x"01d0", -- MOV
    000481 => x"be9e", -- BL
    000482 => x"be4f", -- BL
    000483 => x"3c80", -- SFT
    000484 => x"be4d", -- BL
    000485 => x"2690", -- ORR
    000486 => x"20d5", -- STUB
    000487 => x"c104", -- LDIL
    000488 => x"3dd0", -- SFT
    000489 => x"be96", -- BL
    000490 => x"c105", -- LDIL
    000491 => x"01d0", -- MOV
    000492 => x"be93", -- BL
    000493 => x"c106", -- LDIL
    000494 => x"be43", -- BL
    000495 => x"0180", -- MOV
    000496 => x"be8f", -- BL
    000497 => x"0121", -- INC
    000498 => x"c010", -- LDIL
    000499 => x"1828", -- CMP
    000500 => x"85fa", -- BNE
    000501 => x"c110", -- LDIL
    000502 => x"2ad5", -- CLR
    000503 => x"be3a", -- BL
    000504 => x"0180", -- MOV
    000505 => x"be86", -- BL
    000506 => x"0121", -- INC
    000507 => x"2400", -- LDUB
    000508 => x"02d1", -- INC
    000509 => x"1858", -- CMP
    000510 => x"85f9", -- BNE
    000511 => x"c001", -- LDIL
    000512 => x"ed0c", -- MCR
    000513 => x"c050", -- LDIL
    000514 => x"c83f", -- LDIH
    000515 => x"ed0a", -- MCR
    000516 => x"c00c", -- LDIL
    000517 => x"c801", -- LDIH
    000518 => x"be73", -- BL
    000519 => x"c524", -- LDIL
    000520 => x"c906", -- LDIH
    000521 => x"be0e", -- BL
    000522 => x"c6a0", -- LDIL
    000523 => x"ca80", -- LDIH
    000524 => x"3450", -- GT
    000525 => x"c52e", -- LDIL
    000526 => x"c907", -- LDIH
    000527 => x"be08", -- BL
    000528 => x"c564", -- LDIL
    000529 => x"c907", -- LDIH
    000530 => x"be05", -- BL
    000531 => x"be1e", -- BL
    000532 => x"2800", -- CLR
    000533 => x"3400", -- GT
    000534 => x"bc9e", -- B
    000535 => x"c5ff", -- LDIL
    000536 => x"0270", -- MOV
    000537 => x"bc03", -- B
    000538 => x"29b3", -- CLR
    000539 => x"0270", -- MOV
    000540 => x"7829", -- LDR
    000541 => x"c080", -- LDIL
    000542 => x"ccff", -- LDIH
    000543 => x"2081", -- AND
    000544 => x"3c98", -- SFTS
    000545 => x"8003", -- BEQ
    000546 => x"be0a", -- BL
    000547 => x"bdf9", -- B
    000548 => x"03c0", -- MOV
    000549 => x"343b", -- TEQ
    000550 => x"f707", -- RBAEQ
    000551 => x"0170", -- MOV
    000552 => x"c08d", -- LDIL
    000553 => x"be03", -- BL
    000554 => x"c08a", -- LDIL
    000555 => x"03a0", -- MOV
    000556 => x"ec22", -- MRC
    000557 => x"dc05", -- STB
    000558 => x"b9fe", -- BTS
    000559 => x"ed18", -- MCR
    000560 => x"3470", -- RET
    000561 => x"ec20", -- MRC
    000562 => x"dc8f", -- STBI
    000563 => x"b9fe", -- BTS
    000564 => x"c800", -- LDIH
    000565 => x"3470", -- RET
    000566 => x"0170", -- MOV
    000567 => x"c200", -- LDIL
    000568 => x"c184", -- LDIL
    000569 => x"bff8", -- BL
    000570 => x"c0c6", -- LDIL
    000571 => x"1809", -- CMP
    000572 => x"9003", -- BMI
    000573 => x"c0a0", -- LDIL
    000574 => x"1001", -- SUB
    000575 => x"c0b0", -- LDIL
    000576 => x"1809", -- CMP
    000577 => x"91f8", -- BMI
    000578 => x"c0c6", -- LDIL
    000579 => x"1818", -- CMP
    000580 => x"91f5", -- BMI
    000581 => x"c0b9", -- LDIL
    000582 => x"1818", -- CMP
    000583 => x"a404", -- BLS
    000584 => x"c0c1", -- LDIL
    000585 => x"1809", -- CMP
    000586 => x"a1ef", -- BHI
    000587 => x"0080", -- MOV
    000588 => x"bfe0", -- BL
    000589 => x"c030", -- LDIL
    000590 => x"1090", -- SUB
    000591 => x"c009", -- LDIL
    000592 => x"1809", -- CMP
    000593 => x"a402", -- BLS
    000594 => x"0497", -- DEC
    000595 => x"3e42", -- SFT
    000596 => x"3e42", -- SFT
    000597 => x"3e42", -- SFT
    000598 => x"3e42", -- SFT
    000599 => x"2641", -- ORR
    000600 => x"05b9", -- DECS
    000601 => x"85e0", -- BNE
    000602 => x"3420", -- RET
    000603 => x"0370", -- MOV
    000604 => x"3d42", -- SFT
    000605 => x"3d22", -- SFT
    000606 => x"3d22", -- SFT
    000607 => x"3d22", -- SFT
    000608 => x"be0f", -- BL
    000609 => x"bfcb", -- BL
    000610 => x"3d40", -- SFT
    000611 => x"be0c", -- BL
    000612 => x"bfc8", -- BL
    000613 => x"3d45", -- SFT
    000614 => x"3d25", -- SFT
    000615 => x"3d25", -- SFT
    000616 => x"3d25", -- SFT
    000617 => x"be06", -- BL
    000618 => x"bfc2", -- BL
    000619 => x"0140", -- MOV
    000620 => x"be03", -- BL
    000621 => x"bfbf", -- BL
    000622 => x"3460", -- RET
    000623 => x"c08f", -- LDIL
    000624 => x"2121", -- AND
    000625 => x"c089", -- LDIL
    000626 => x"181a", -- CMP
    000627 => x"8803", -- BCS
    000628 => x"c0b0", -- LDIL
    000629 => x"bc02", -- B
    000630 => x"c0b7", -- LDIL
    000631 => x"0892", -- ADD
    000632 => x"3470", -- RET
    000633 => x"ed0b", -- MCR
    000634 => x"ec22", -- MRC
    000635 => x"dc03", -- STB
    000636 => x"b9fe", -- BTS
    000637 => x"ec23", -- MRC
    000638 => x"3470", -- RET
    000639 => x"00f0", -- MOV
    000640 => x"c050", -- LDIL
    000641 => x"c837", -- LDIH
    000642 => x"ed0a", -- MCR
    000643 => x"c001", -- LDIL
    000644 => x"ed0c", -- MCR
    000645 => x"c006", -- LDIL
    000646 => x"bff3", -- BL
    000647 => x"c050", -- LDIL
    000648 => x"c83f", -- LDIH
    000649 => x"ed0a", -- MCR
    000650 => x"c000", -- LDIL
    000651 => x"c805", -- LDIH
    000652 => x"bfed", -- BL
    000653 => x"dc01", -- STB
    000654 => x"b80a", -- BTS
    000655 => x"c554", -- LDIL
    000656 => x"c907", -- LDIH
    000657 => x"bf86", -- BL
    000658 => x"c564", -- LDIL
    000659 => x"c907", -- LDIH
    000660 => x"bf83", -- BL
    000661 => x"bf9c", -- BL
    000662 => x"2800", -- CLR
    000663 => x"3400", -- GT
    000664 => x"c040", -- LDIL
    000665 => x"c83f", -- LDIH
    000666 => x"ed0a", -- MCR
    000667 => x"c001", -- LDIL
    000668 => x"ed0c", -- MCR
    000669 => x"3c20", -- SFT
    000670 => x"c802", -- LDIH
    000671 => x"bfda", -- BL
    000672 => x"03a0", -- MOV
    000673 => x"cb80", -- LDIH
    000674 => x"3ff0", -- SFT
    000675 => x"0030", -- MOV
    000676 => x"c800", -- LDIH
    000677 => x"2407", -- ORR
    000678 => x"bfd3", -- BL
    000679 => x"2800", -- CLR
    000680 => x"ed0c", -- MCR
    000681 => x"c050", -- LDIL
    000682 => x"c83f", -- LDIH
    000683 => x"ed0a", -- MCR
    000684 => x"c001", -- LDIL
    000685 => x"ed0c", -- MCR
    000686 => x"c000", -- LDIL
    000687 => x"c805", -- LDIH
    000688 => x"bfc9", -- BL
    000689 => x"dc00", -- STB
    000690 => x"b9fc", -- BTS
    000691 => x"3410", -- RET
    000692 => x"00f0", -- MOV
    000693 => x"c040", -- LDIL
    000694 => x"c83f", -- LDIH
    000695 => x"ed0a", -- MCR
    000696 => x"c001", -- LDIL
    000697 => x"ed0c", -- MCR
    000698 => x"3c20", -- SFT
    000699 => x"c803", -- LDIH
    000700 => x"bfbd", -- BL
    000701 => x"0020", -- MOV
    000702 => x"c800", -- LDIH
    000703 => x"3c00", -- SFT
    000704 => x"bfb9", -- BL
    000705 => x"29b3", -- CLR
    000706 => x"ed3c", -- MCR
    000707 => x"0180", -- MOV
    000708 => x"c980", -- LDIH
    000709 => x"3410", -- RET
    000710 => x"c54e", -- LDIL
    000711 => x"c906", -- LDIH
    000712 => x"bf52", -- BL
    000713 => x"bf6d", -- BL
    000714 => x"edca", -- MCR
    000715 => x"bf6b", -- BL
    000716 => x"edc9", -- MCR
    000717 => x"bf64", -- BL
    000718 => x"c08d", -- LDIL
    000719 => x"1809", -- CMP
    000720 => x"8005", -- BEQ
    000721 => x"c088", -- LDIL
    000722 => x"1809", -- CMP
    000723 => x"8009", -- BEQ
    000724 => x"bdf9", -- B
    000725 => x"be0b", -- BL
    000726 => x"0300", -- MOV
    000727 => x"c572", -- LDIL
    000728 => x"c906", -- LDIH
    000729 => x"bf41", -- BL
    000730 => x"0260", -- MOV
    000731 => x"bf80", -- BL
    000732 => x"bf4b", -- BL
    000733 => x"c6c6", -- LDIL
    000734 => x"ca80", -- LDIH
    000735 => x"3450", -- GT
    000736 => x"e5b0", -- CDP
    000737 => x"ec30", -- MRC
    000738 => x"dc06", -- STB
    000739 => x"b9fe", -- BTS
    000740 => x"ec34", -- MRC
    000741 => x"3470", -- RET
    000742 => x"4174", -- .DW
    000743 => x"6c61", -- .DW
    000744 => x"732d", -- .DW
    000745 => x"324b", -- .DW
    000746 => x"2042", -- .DW
    000747 => x"6f6f", -- .DW
    000748 => x"746c", -- .DW
    000749 => x"6f61", -- .DW
    000750 => x"6465", -- .DW
    000751 => x"7220", -- .DW
    000752 => x"2d20", -- .DW
    000753 => x"5632", -- .DW
    000754 => x"3031", -- .DW
    000755 => x"3430", -- .DW
    000756 => x"3431", -- .DW
    000757 => x"300d", -- .DW
    000758 => x"0a62", -- .DW
    000759 => x"7920", -- .DW
    000760 => x"5374", -- .DW
    000761 => x"6570", -- .DW
    000762 => x"6861", -- .DW
    000763 => x"6e20", -- .DW
    000764 => x"4e6f", -- .DW
    000765 => x"6c74", -- .DW
    000766 => x"696e", -- .DW
    000767 => x"672c", -- .DW
    000768 => x"2073", -- .DW
    000769 => x"746e", -- .DW
    000770 => x"6f6c", -- .DW
    000771 => x"7469", -- .DW
    000772 => x"6e67", -- .DW
    000773 => x"4067", -- .DW
    000774 => x"6d61", -- .DW
    000775 => x"696c", -- .DW
    000776 => x"2e63", -- .DW
    000777 => x"6f6d", -- .DW
    000778 => x"0d0a", -- .DW
    000779 => x"7777", -- .DW
    000780 => x"772e", -- .DW
    000781 => x"6f70", -- .DW
    000782 => x"656e", -- .DW
    000783 => x"636f", -- .DW
    000784 => x"7265", -- .DW
    000785 => x"732e", -- .DW
    000786 => x"6f72", -- .DW
    000787 => x"672f", -- .DW
    000788 => x"7072", -- .DW
    000789 => x"6f6a", -- .DW
    000790 => x"6563", -- .DW
    000791 => x"742c", -- .DW
    000792 => x"6174", -- .DW
    000793 => x"6c61", -- .DW
    000794 => x"735f", -- .DW
    000795 => x"636f", -- .DW
    000796 => x"7265", -- .DW
    000797 => x"0d0a", -- .DW
    000798 => x"0000", -- .DW
    000799 => x"426f", -- .DW
    000800 => x"6f74", -- .DW
    000801 => x"6c6f", -- .DW
    000802 => x"6164", -- .DW
    000803 => x"6572", -- .DW
    000804 => x"2040", -- .DW
    000805 => x"2030", -- .DW
    000806 => x"7800", -- .DW
    000807 => x"436c", -- .DW
    000808 => x"6f63", -- .DW
    000809 => x"6b20", -- .DW
    000810 => x"2848", -- .DW
    000811 => x"7a29", -- .DW
    000812 => x"3a20", -- .DW
    000813 => x"3078", -- .DW
    000814 => x"0000", -- .DW
    000815 => x"426f", -- .DW
    000816 => x"6f74", -- .DW
    000817 => x"696e", -- .DW
    000818 => x"672e", -- .DW
    000819 => x"2e2e", -- .DW
    000820 => x"0000", -- .DW
    000821 => x"4275", -- .DW
    000822 => x"726e", -- .DW
    000823 => x"696e", -- .DW
    000824 => x"6720", -- .DW
    000825 => x"4545", -- .DW
    000826 => x"5052", -- .DW
    000827 => x"4f4d", -- .DW
    000828 => x"0000", -- .DW
    000829 => x"5761", -- .DW
    000830 => x"6974", -- .DW
    000831 => x"696e", -- .DW
    000832 => x"6720", -- .DW
    000833 => x"666f", -- .DW
    000834 => x"7220", -- .DW
    000835 => x"696d", -- .DW
    000836 => x"6167", -- .DW
    000837 => x"6520", -- .DW
    000838 => x"6461", -- .DW
    000839 => x"7461", -- .DW
    000840 => x"2e2e", -- .DW
    000841 => x"2e00", -- .DW
    000842 => x"5374", -- .DW
    000843 => x"6172", -- .DW
    000844 => x"7469", -- .DW
    000845 => x"6e67", -- .DW
    000846 => x"2069", -- .DW
    000847 => x"6d61", -- .DW
    000848 => x"6765", -- .DW
    000849 => x"2000", -- .DW
    000850 => x"446f", -- .DW
    000851 => x"776e", -- .DW
    000852 => x"6c6f", -- .DW
    000853 => x"6164", -- .DW
    000854 => x"2063", -- .DW
    000855 => x"6f6d", -- .DW
    000856 => x"706c", -- .DW
    000857 => x"6574", -- .DW
    000858 => x"6564", -- .DW
    000859 => x"2100", -- .DW
    000860 => x"456e", -- .DW
    000861 => x"7465", -- .DW
    000862 => x"7220", -- .DW
    000863 => x"7061", -- .DW
    000864 => x"6765", -- .DW
    000865 => x"2028", -- .DW
    000866 => x"3468", -- .DW
    000867 => x"6578", -- .DW
    000868 => x"293a", -- .DW
    000869 => x"2030", -- .DW
    000870 => x"7800", -- .DW
    000871 => x"456e", -- .DW
    000872 => x"7465", -- .DW
    000873 => x"7220", -- .DW
    000874 => x"6164", -- .DW
    000875 => x"6472", -- .DW
    000876 => x"2028", -- .DW
    000877 => x"3868", -- .DW
    000878 => x"6578", -- .DW
    000879 => x"293a", -- .DW
    000880 => x"2030", -- .DW
    000881 => x"7800", -- .DW
    000882 => x"4368", -- .DW
    000883 => x"6563", -- .DW
    000884 => x"6b73", -- .DW
    000885 => x"756d", -- .DW
    000886 => x"3a20", -- .DW
    000887 => x"3078", -- .DW
    000888 => x"0000", -- .DW
    000889 => x"0d0a", -- .DW
    000890 => x"2d3e", -- .DW
    000891 => x"2030", -- .DW
    000892 => x"7800", -- .DW
    000893 => x"636d", -- .DW
    000894 => x"642f", -- .DW
    000895 => x"626f", -- .DW
    000896 => x"6f74", -- .DW
    000897 => x"2d73", -- .DW
    000898 => x"7769", -- .DW
    000899 => x"7463", -- .DW
    000900 => x"6800", -- .DW
    000901 => x"2030", -- .DW
    000902 => x"2f27", -- .DW
    000903 => x"3030", -- .DW
    000904 => x"273a", -- .DW
    000905 => x"2052", -- .DW
    000906 => x"6573", -- .DW
    000907 => x"7461", -- .DW
    000908 => x"7274", -- .DW
    000909 => x"2063", -- .DW
    000910 => x"6f6e", -- .DW
    000911 => x"736f", -- .DW
    000912 => x"6c65", -- .DW
    000913 => x"0d0a", -- .DW
    000914 => x"2031", -- .DW
    000915 => x"2f27", -- .DW
    000916 => x"3031", -- .DW
    000917 => x"273a", -- .DW
    000918 => x"2042", -- .DW
    000919 => x"6f6f", -- .DW
    000920 => x"7420", -- .DW
    000921 => x"6672", -- .DW
    000922 => x"6f6d", -- .DW
    000923 => x"2055", -- .DW
    000924 => x"4152", -- .DW
    000925 => x"540d", -- .DW
    000926 => x"0a20", -- .DW
    000927 => x"322f", -- .DW
    000928 => x"2731", -- .DW
    000929 => x"3027", -- .DW
    000930 => x"3a20", -- .DW
    000931 => x"426f", -- .DW
    000932 => x"6f74", -- .DW
    000933 => x"2066", -- .DW
    000934 => x"726f", -- .DW
    000935 => x"6d20", -- .DW
    000936 => x"4545", -- .DW
    000937 => x"5052", -- .DW
    000938 => x"4f4d", -- .DW
    000939 => x"0d0a", -- .DW
    000940 => x"2033", -- .DW
    000941 => x"2f27", -- .DW
    000942 => x"3131", -- .DW
    000943 => x"273a", -- .DW
    000944 => x"2042", -- .DW
    000945 => x"6f6f", -- .DW
    000946 => x"7420", -- .DW
    000947 => x"6672", -- .DW
    000948 => x"6f6d", -- .DW
    000949 => x"206d", -- .DW
    000950 => x"656d", -- .DW
    000951 => x"6f72", -- .DW
    000952 => x"7900", -- .DW
    000953 => x"2070", -- .DW
    000954 => x"3a20", -- .DW
    000955 => x"4275", -- .DW
    000956 => x"726e", -- .DW
    000957 => x"2045", -- .DW
    000958 => x"4550", -- .DW
    000959 => x"524f", -- .DW
    000960 => x"4d00", -- .DW
    000961 => x"2064", -- .DW
    000962 => x"3a20", -- .DW
    000963 => x"5241", -- .DW
    000964 => x"4d20", -- .DW
    000965 => x"6475", -- .DW
    000966 => x"6d70", -- .DW
    000967 => x"0000", -- .DW
    000968 => x"2072", -- .DW
    000969 => x"3a20", -- .DW
    000970 => x"5265", -- .DW
    000971 => x"7365", -- .DW
    000972 => x"7400", -- .DW
    000973 => x"2077", -- .DW
    000974 => x"3a20", -- .DW
    000975 => x"5742", -- .DW
    000976 => x"2064", -- .DW
    000977 => x"756d", -- .DW
    000978 => x"7000", -- .DW
    000979 => x"636d", -- .DW
    000980 => x"643a", -- .DW
    000981 => x"3e20", -- .DW
    000982 => x"0000", -- .DW
    000983 => x"494d", -- .DW
    000984 => x"4147", -- .DW
    000985 => x"4520", -- .DW
    000986 => x"4552", -- .DW
    000987 => x"5221", -- .DW
    000988 => x"0000", -- .DW
    000989 => x"0d0a", -- .DW
    000990 => x"4952", -- .DW
    000991 => x"5120", -- .DW
    000992 => x"4552", -- .DW
    000993 => x"5221", -- .DW
    000994 => x"0000", -- .DW
    000995 => x"4348", -- .DW
    000996 => x"4543", -- .DW
    000997 => x"4b53", -- .DW
    000998 => x"554d", -- .DW
    000999 => x"2045", -- .DW
    001000 => x"5252", -- .DW
    001001 => x"2100", -- .DW
    001002 => x"5350", -- .DW
    001003 => x"492f", -- .DW
    001004 => x"4545", -- .DW
    001005 => x"5052", -- .DW
    001006 => x"4f4d", -- .DW
    001007 => x"2045", -- .DW
    001008 => x"5252", -- .DW
    001009 => x"2100", -- .DW
    001010 => x"5072", -- .DW
    001011 => x"6573", -- .DW
    001012 => x"7320", -- .DW
    001013 => x"616e", -- .DW
    001014 => x"7920", -- .DW
    001015 => x"6b65", -- .DW
    001016 => x"7900", -- .DW
    others => x"0000"  -- NOP
	);
	------------------------------------------------------

begin

	-- Memory Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		MEM_FILE_ACCESS: process(CLK_I)
		begin
			if rising_edge(CLK_I) then
				-- Data Read --
				if (D_EN_I = '1') then -- valid access
					if (word_mode_en_c = true) then -- read data access
						D_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(D_ADR_I(log2_mem_size_c-1 downto 0))));
					else
						D_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(D_ADR_I(log2_mem_size_c downto 1))));
					end if;
				end if;
				-- Instruction Read --
				if (I_EN_I = '1') then
					if (word_mode_en_c = true) then
						I_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(I_ADR_I(log2_mem_size_c-1 downto 0))));
					else
						I_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(I_ADR_I(log2_mem_size_c downto 1))));
					end if;
				end if;
			end if;
		end process MEM_FILE_ACCESS;



end BOOT_MEM_STRUCTURE;
