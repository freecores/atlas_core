000000 => x"bc0b", -- B
000001 => x"bc04", -- B
000002 => x"bc03", -- B
000003 => x"bc02", -- B
000004 => x"bc01", -- B
000005 => x"be31", -- BL
000006 => x"c110", -- LDIL
000007 => x"c901", -- LDIH
000008 => x"be21", -- BL
000009 => x"be2d", -- BL
000010 => x"bc00", -- B
000011 => x"c12c", -- LDIL
000012 => x"c901", -- LDIH
000013 => x"be19", -- BL
000014 => x"c144", -- LDIL
000015 => x"c901", -- LDIH
000016 => x"be19", -- BL
000017 => x"be34", -- BL
000018 => x"ec4d", -- MCR
000019 => x"be23", -- BL
000020 => x"c160", -- LDIL
000021 => x"c901", -- LDIH
000022 => x"be13", -- BL
000023 => x"be2e", -- BL
000024 => x"d24f", -- CBR
000025 => x"ec4e", -- MCR
000026 => x"be1c", -- BL
000027 => x"c0b0", -- LDIL
000028 => x"be1f", -- BL
000029 => x"c0f8", -- LDIL
000030 => x"be1d", -- BL
000031 => x"ee05", -- MRC
000032 => x"be4a", -- BL
000033 => x"be15", -- BL
000034 => x"ec20", -- MRC
000035 => x"dc0f", -- STB
000036 => x"b9ea", -- BTS
000037 => x"bdf6", -- B
000038 => x"c5ff", -- LDIL
000039 => x"0270", -- MOV
000040 => x"bc03", -- B
000041 => x"29b3", -- CLR
000042 => x"0270", -- MOV
000043 => x"7829", -- LDR
000044 => x"c080", -- LDIL
000045 => x"ccff", -- LDIH
000046 => x"2081", -- AND
000047 => x"3c98", -- SFTS
000048 => x"8003", -- BEQ
000049 => x"be0a", -- BL
000050 => x"bdf9", -- B
000051 => x"03c0", -- MOV
000052 => x"343b", -- TEQ
000053 => x"f707", -- RBAEQ
000054 => x"0170", -- MOV
000055 => x"c08d", -- LDIL
000056 => x"be03", -- BL
000057 => x"c08a", -- LDIL
000058 => x"03a0", -- MOV
000059 => x"ec22", -- MRC
000060 => x"dc05", -- STB
000061 => x"b9fe", -- BTS
000062 => x"ed18", -- MCR
000063 => x"3470", -- RET
000064 => x"ec20", -- MRC
000065 => x"dc8f", -- STBI
000066 => x"b9fe", -- BTS
000067 => x"c800", -- LDIH
000068 => x"3470", -- RET
000069 => x"0170", -- MOV
000070 => x"c200", -- LDIL
000071 => x"c184", -- LDIL
000072 => x"bff8", -- BL
000073 => x"c0c6", -- LDIL
000074 => x"1809", -- CMP
000075 => x"9003", -- BMI
000076 => x"c0a0", -- LDIL
000077 => x"1001", -- SUB
000078 => x"c0b0", -- LDIL
000079 => x"1809", -- CMP
000080 => x"91f8", -- BMI
000081 => x"c0c6", -- LDIL
000082 => x"1818", -- CMP
000083 => x"91f5", -- BMI
000084 => x"c0b9", -- LDIL
000085 => x"1818", -- CMP
000086 => x"a404", -- BLS
000087 => x"c0c1", -- LDIL
000088 => x"1809", -- CMP
000089 => x"a1ef", -- BHI
000090 => x"0080", -- MOV
000091 => x"bfe0", -- BL
000092 => x"c030", -- LDIL
000093 => x"1090", -- SUB
000094 => x"c009", -- LDIL
000095 => x"1809", -- CMP
000096 => x"a402", -- BLS
000097 => x"0497", -- DEC
000098 => x"3e42", -- SFT
000099 => x"3e42", -- SFT
000100 => x"3e42", -- SFT
000101 => x"3e42", -- SFT
000102 => x"2641", -- ORR
000103 => x"05b9", -- DECS
000104 => x"85e0", -- BNE
000105 => x"3420", -- RET
000106 => x"0370", -- MOV
000107 => x"3d42", -- SFT
000108 => x"3d22", -- SFT
000109 => x"3d22", -- SFT
000110 => x"3d22", -- SFT
000111 => x"be0f", -- BL
000112 => x"bfcb", -- BL
000113 => x"3d40", -- SFT
000114 => x"be0c", -- BL
000115 => x"bfc8", -- BL
000116 => x"3d45", -- SFT
000117 => x"3d25", -- SFT
000118 => x"3d25", -- SFT
000119 => x"3d25", -- SFT
000120 => x"be06", -- BL
000121 => x"bfc2", -- BL
000122 => x"0140", -- MOV
000123 => x"be03", -- BL
000124 => x"bfbf", -- BL
000125 => x"3460", -- RET
000126 => x"c08f", -- LDIL
000127 => x"2121", -- AND
000128 => x"c089", -- LDIL
000129 => x"181a", -- CMP
000130 => x"8803", -- BCS
000131 => x"c0b0", -- LDIL
000132 => x"bc02", -- B
000133 => x"c0b7", -- LDIL
000134 => x"0892", -- ADD
000135 => x"3470", -- RET
000136 => x"4578", -- .DW
000137 => x"6365", -- .DW
000138 => x"7074", -- .DW
000139 => x"696f", -- .DW
000140 => x"6e2f", -- .DW
000141 => x"696e", -- .DW
000142 => x"7465", -- .DW
000143 => x"7272", -- .DW
000144 => x"7570", -- .DW
000145 => x"7420", -- .DW
000146 => x"6572", -- .DW
000147 => x"726f", -- .DW
000148 => x"7221", -- .DW
000149 => x"0000", -- .DW
000150 => x"5261", -- .DW
000151 => x"6e64", -- .DW
000152 => x"6f6d", -- .DW
000153 => x"204e", -- .DW
000154 => x"756d", -- .DW
000155 => x"6265", -- .DW
000156 => x"7220", -- .DW
000157 => x"4765", -- .DW
000158 => x"6e65", -- .DW
000159 => x"7261", -- .DW
000160 => x"746f", -- .DW
000161 => x"7200", -- .DW
000162 => x"456e", -- .DW
000163 => x"7465", -- .DW
000164 => x"7220", -- .DW
000165 => x"4c46", -- .DW
000166 => x"5352", -- .DW
000167 => x"2073", -- .DW
000168 => x"6565", -- .DW
000169 => x"6420", -- .DW
000170 => x"2834", -- .DW
000171 => x"6865", -- .DW
000172 => x"7829", -- .DW
000173 => x"3a20", -- .DW
000174 => x"3078", -- .DW
000175 => x"0000", -- .DW
000176 => x"456e", -- .DW
000177 => x"7465", -- .DW
000178 => x"7220", -- .DW
000179 => x"4c46", -- .DW
000180 => x"5352", -- .DW
000181 => x"2074", -- .DW
000182 => x"6170", -- .DW
000183 => x"7320", -- .DW
000184 => x"2834", -- .DW
000185 => x"6865", -- .DW
000186 => x"7829", -- .DW
000187 => x"3a20", -- .DW
000188 => x"3078", -- .DW
000189 => x"0000", -- .DW
others => x"0000"  -- NOP