-- ########################################################
-- #         << ATLAS Project - Bootloader ROM >>         #
-- # **************************************************** #
-- #  Initialized with boot loader.                       #
-- # **************************************************** #
-- #  Last modified: 08.03.2014                           #
-- # **************************************************** #
-- #  by Stephan Nolting 4788, Hanover, Germany           #
-- ########################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.atlas_core_package.all;

entity BOOT_MEM is
	port	(
				-- Host Interface --
				CLK_I           : in  std_logic; -- global clock line
				I_ADR_I         : in  std_logic_vector(15 downto 0); -- instruction adr
				I_EN_I          : in  std_logic; -- IR update
				I_DAT_O         : out std_logic_vector(15 downto 0); -- instruction out
				D_EN_I          : in  std_logic; -- access enable
				D_RW_I          : in  std_logic; -- read/write
				D_ADR_I         : in  std_logic_vector(15 downto 0); -- data adr
				D_DAT_I         : in  std_logic_vector(15 downto 0); -- data in
				D_DAT_O         : out std_logic_vector(15 downto 0)  -- data out
			);
end BOOT_MEM;

architecture BOOT_MEM_STRUCTURE of BOOT_MEM is

	-- Internal constants(configuration --
	constant mem_size_c      : natural := 2048; -- 2kB
	constant log2_mem_size_c : natural := log2(mem_size_c/2); -- address width (word boundary!)

	-- Memory Type --
	type mem_file_t is array (0 to (mem_size_c/2)-1) of std_logic_vector(15 downto 0); -- word mem!

	-- MEMORY IMAGE (Bootloader Program) --
	------------------------------------------------------
	constant BOOT_MEM_FILE_C : mem_file_t :=
	(
		000000 => x"bc0e", -- B
		000001 => x"bc04", -- B
		000002 => x"bc03", -- B
		000003 => x"bc02", -- B
		000004 => x"bc01", -- B
		000005 => x"c000", -- LDIL
		000006 => x"cc00", -- LDIH
		000007 => x"ec8a", -- MCR
		000008 => x"ed0f", -- MCR
		000009 => x"be8f", -- BL
		000010 => x"c524", -- LDIL
		000011 => x"c907", -- LDIH
		000012 => x"be8a", -- BL
		000013 => x"bc00", -- B
		000014 => x"c000", -- LDIL
		000015 => x"cc78", -- LDIH
		000016 => x"1c00", -- STSR
		000017 => x"ec11", -- MRC
		000018 => x"ec88", -- MCR
		000019 => x"ec8a", -- MCR
		000020 => x"c000", -- LDIL
		000021 => x"ec08", -- MCR
		000022 => x"ec09", -- MCR
		000023 => x"ec0a", -- MCR
		000024 => x"ec0b", -- MCR
		000025 => x"ec0c", -- MCR
		000026 => x"ec0d", -- MCR
		000027 => x"ec0e", -- MCR
		000028 => x"ec00", -- MRC
		000029 => x"c801", -- LDIH
		000030 => x"ed0f", -- MCR
		000031 => x"ec17", -- MRC
		000032 => x"ec97", -- MRC
		000033 => x"c160", -- LDIL
		000034 => x"c909", -- LDIH
		000035 => x"c18f", -- LDIL
		000036 => x"0923", -- ADD
		000037 => x"29b3", -- CLR
		000038 => x"2a44", -- CLR
		000039 => x"100a", -- SUBS
		000040 => x"149b", -- SBCS
		000041 => x"9003", -- BMI
		000042 => x"0241", -- INC
		000043 => x"bdfc", -- B
		000044 => x"ed49", -- MCR
		000045 => x"ec22", -- MRC
		000046 => x"d406", -- SBR
		000047 => x"ed0a", -- MCR
		000048 => x"be68", -- BL
		000049 => x"be67", -- BL
		000050 => x"c510", -- LDIL
		000051 => x"c905", -- LDIH
		000052 => x"be62", -- BL
		000053 => x"c53a", -- LDIL
		000054 => x"c905", -- LDIH
		000055 => x"be5f", -- BL
		000056 => x"c562", -- LDIL
		000057 => x"c905", -- LDIH
		000058 => x"be5c", -- BL
		000059 => x"be5d", -- BL
		000060 => x"c108", -- LDIL
		000061 => x"c906", -- LDIH
		000062 => x"be59", -- BL
		000063 => x"ee11", -- MRC
		000064 => x"be5b", -- BL
		000065 => x"be57", -- BL
		000066 => x"c11e", -- LDIL
		000067 => x"c906", -- LDIH
		000068 => x"be53", -- BL
		000069 => x"ee97", -- MRC
		000070 => x"ee17", -- MRC
		000071 => x"be54", -- BL
		000072 => x"0250", -- MOV
		000073 => x"be52", -- BL
		000074 => x"be4e", -- BL
		000075 => x"ec27", -- MRC
		000076 => x"c083", -- LDIL
		000077 => x"2001", -- AND
		000078 => x"c330", -- LDIL
		000079 => x"0b60", -- ADD
		000080 => x"bc22", -- B
		000081 => x"be47", -- BL
		000082 => x"c568", -- LDIL
		000083 => x"c906", -- LDIH
		000084 => x"be42", -- BL
		000085 => x"c57c", -- LDIL
		000086 => x"c906", -- LDIH
		000087 => x"be3f", -- BL
		000088 => x"c116", -- LDIL
		000089 => x"c907", -- LDIH
		000090 => x"be3c", -- BL
		000091 => x"c12e", -- LDIL
		000092 => x"c907", -- LDIH
		000093 => x"be39", -- BL
		000094 => x"c148", -- LDIL
		000095 => x"c907", -- LDIH
		000096 => x"be36", -- BL
		000097 => x"c162", -- LDIL
		000098 => x"c907", -- LDIH
		000099 => x"be33", -- BL
		000100 => x"c176", -- LDIL
		000101 => x"c907", -- LDIH
		000102 => x"be30", -- BL
		000103 => x"c504", -- LDIL
		000104 => x"c907", -- LDIH
		000105 => x"be2d", -- BL
		000106 => x"c50e", -- LDIL
		000107 => x"c907", -- LDIH
		000108 => x"be2b", -- BL
		000109 => x"be2d", -- BL
		000110 => x"0300", -- MOV
		000111 => x"00e0", -- MOV
		000112 => x"be29", -- BL
		000113 => x"be27", -- BL
		000114 => x"c0b0", -- LDIL
		000115 => x"181e", -- CMP
		000116 => x"81dd", -- BEQ
		000117 => x"c0b1", -- LDIL
		000118 => x"181e", -- CMP
		000119 => x"8076", -- BEQ
		000120 => x"c0b2", -- LDIL
		000121 => x"181e", -- CMP
		000122 => x"8022", -- BEQ
		000123 => x"c0b3", -- LDIL
		000124 => x"181e", -- CMP
		000125 => x"8013", -- BEQ
		000126 => x"c2f8", -- LDIL
		000127 => x"ca83", -- LDIH
		000128 => x"c0f0", -- LDIL
		000129 => x"181e", -- CMP
		000130 => x"f705", -- RBAEQ
		000131 => x"c6f6", -- LDIL
		000132 => x"ca82", -- LDIH
		000133 => x"c0e4", -- LDIL
		000134 => x"181e", -- CMP
		000135 => x"f705", -- RBAEQ
		000136 => x"c0f2", -- LDIL
		000137 => x"181e", -- CMP
		000138 => x"85e0", -- BNE
		000139 => x"2800", -- CLR
		000140 => x"c080", -- LDIL
		000141 => x"cc80", -- LDIH
		000142 => x"ec99", -- MCR
		000143 => x"3400", -- GT
		000144 => x"c508", -- LDIL
		000145 => x"c906", -- LDIH
		000146 => x"be04", -- BL
		000147 => x"2800", -- CLR
		000148 => x"2100", -- STUB
		000149 => x"bcb1", -- B
		000150 => x"bca7", -- B
		000151 => x"bca7", -- B
		000152 => x"bca7", -- B
		000153 => x"bca7", -- B
		000154 => x"bca7", -- B
		000155 => x"bcaa", -- B
		000156 => x"c134", -- LDIL
		000157 => x"c906", -- LDIH
		000158 => x"be9f", -- BL
		000159 => x"c100", -- LDIL
		000160 => x"bea2", -- BL
		000161 => x"3eb0", -- SFT
		000162 => x"c101", -- LDIL
		000163 => x"be9f", -- BL
		000164 => x"26d3", -- ORR
		000165 => x"c47e", -- LDIL
		000166 => x"cc4a", -- LDIH
		000167 => x"180d", -- CMP
		000168 => x"849b", -- BNE
		000169 => x"c102", -- LDIL
		000170 => x"be98", -- BL
		000171 => x"3eb0", -- SFT
		000172 => x"c103", -- LDIL
		000173 => x"be95", -- BL
		000174 => x"26d3", -- ORR
		000175 => x"2055", -- STUB
		000176 => x"c104", -- LDIL
		000177 => x"be91", -- BL
		000178 => x"3eb0", -- SFT
		000179 => x"c105", -- LDIL
		000180 => x"be8e", -- BL
		000181 => x"26d3", -- ORR
		000182 => x"20d5", -- STUB
		000183 => x"c106", -- LDIL
		000184 => x"be8a", -- BL
		000185 => x"3eb0", -- SFT
		000186 => x"c107", -- LDIL
		000187 => x"be87", -- BL
		000188 => x"26d3", -- ORR
		000189 => x"2155", -- STUB
		000190 => x"c108", -- LDIL
		000191 => x"be83", -- BL
		000192 => x"3eb0", -- SFT
		000193 => x"c109", -- LDIL
		000194 => x"be80", -- BL
		000195 => x"26d3", -- ORR
		000196 => x"21d5", -- STUB
		000197 => x"c10a", -- LDIL
		000198 => x"be7c", -- BL
		000199 => x"3eb0", -- SFT
		000200 => x"c10b", -- LDIL
		000201 => x"be79", -- BL
		000202 => x"26d3", -- ORR
		000203 => x"2255", -- STUB
		000204 => x"c10c", -- LDIL
		000205 => x"be75", -- BL
		000206 => x"3eb0", -- SFT
		000207 => x"c10d", -- LDIL
		000208 => x"be72", -- BL
		000209 => x"26d3", -- ORR
		000210 => x"22d5", -- STUB
		000211 => x"c10e", -- LDIL
		000212 => x"be6e", -- BL
		000213 => x"3eb0", -- SFT
		000214 => x"c10f", -- LDIL
		000215 => x"be6b", -- BL
		000216 => x"26d3", -- ORR
		000217 => x"2355", -- STUB
		000218 => x"c300", -- LDIL
		000219 => x"ecea", -- MCR
		000220 => x"23e6", -- STUB
		000221 => x"c010", -- LDIL
		000222 => x"0960", -- ADD
		000223 => x"be63", -- BL
		000224 => x"3eb0", -- SFT
		000225 => x"c011", -- LDIL
		000226 => x"0960", -- ADD
		000227 => x"be5f", -- BL
		000228 => x"26d3", -- ORR
		000229 => x"7eea", -- STR
		000230 => x"2477", -- LDUB
		000231 => x"2805", -- EOR
		000232 => x"2380", -- STUB
		000233 => x"2400", -- LDUB
		000234 => x"1868", -- CMP
		000235 => x"85f2", -- BNE
		000236 => x"bc41", -- B
		000237 => x"c14c", -- LDIL
		000238 => x"c906", -- LDIH
		000239 => x"be4e", -- BL
		000240 => x"c16e", -- LDIL
		000241 => x"c906", -- LDIH
		000242 => x"be4b", -- BL
		000243 => x"be4e", -- BL
		000244 => x"3c80", -- SFT
		000245 => x"be4c", -- BL
		000246 => x"2490", -- ORR
		000247 => x"c47e", -- LDIL
		000248 => x"cc4a", -- LDIH
		000249 => x"1818", -- CMP
		000250 => x"8449", -- BNE
		000251 => x"be46", -- BL
		000252 => x"3c80", -- SFT
		000253 => x"be44", -- BL
		000254 => x"2490", -- ORR
		000255 => x"3c94", -- SFT
		000256 => x"2011", -- STUB
		000257 => x"be40", -- BL
		000258 => x"3c80", -- SFT
		000259 => x"be3e", -- BL
		000260 => x"2490", -- ORR
		000261 => x"2091", -- STUB
		000262 => x"be3b", -- BL
		000263 => x"3c80", -- SFT
		000264 => x"be39", -- BL
		000265 => x"2490", -- ORR
		000266 => x"2111", -- STUB
		000267 => x"be36", -- BL
		000268 => x"3c80", -- SFT
		000269 => x"be34", -- BL
		000270 => x"2490", -- ORR
		000271 => x"2191", -- STUB
		000272 => x"be31", -- BL
		000273 => x"3c80", -- SFT
		000274 => x"be2f", -- BL
		000275 => x"2490", -- ORR
		000276 => x"2211", -- STUB
		000277 => x"be2c", -- BL
		000278 => x"3c80", -- SFT
		000279 => x"be2a", -- BL
		000280 => x"2490", -- ORR
		000281 => x"2291", -- STUB
		000282 => x"be27", -- BL
		000283 => x"3c80", -- SFT
		000284 => x"be25", -- BL
		000285 => x"2490", -- ORR
		000286 => x"2311", -- STUB
		000287 => x"2ad5", -- CLR
		000288 => x"ecda", -- MCR
		000289 => x"23d5", -- STUB
		000290 => x"be1f", -- BL
		000291 => x"3c80", -- SFT
		000292 => x"be1d", -- BL
		000293 => x"2490", -- ORR
		000294 => x"7cda", -- STR
		000295 => x"2477", -- LDUB
		000296 => x"2801", -- EOR
		000297 => x"2380", -- STUB
		000298 => x"2400", -- LDUB
		000299 => x"1858", -- CMP
		000300 => x"85f6", -- BNE
		000301 => x"c000", -- LDIL
		000302 => x"cc00", -- LDIH
		000303 => x"ec8a", -- MCR
		000304 => x"2477", -- LDUB
		000305 => x"2491", -- LDUB
		000306 => x"1809", -- CMP
		000307 => x"8013", -- BEQ
		000308 => x"c530", -- LDIL
		000309 => x"c907", -- LDIH
		000310 => x"be07", -- BL
		000311 => x"c552", -- LDIL
		000312 => x"c907", -- LDIH
		000313 => x"be04", -- BL
		000314 => x"be07", -- BL
		000315 => x"2800", -- CLR
		000316 => x"3400", -- GT
		000317 => x"bcdc", -- B
		000318 => x"bcde", -- B
		000319 => x"bcea", -- B
		000320 => x"bcee", -- B
		000321 => x"bcf2", -- B
		000322 => x"bc78", -- B
		000323 => x"bccc", -- B
		000324 => x"bd26", -- B
		000325 => x"bc76", -- B
		000326 => x"c520", -- LDIL
		000327 => x"c906", -- LDIH
		000328 => x"bed4", -- BL
		000329 => x"24aa", -- LDUBS
		000330 => x"8024", -- BEQ
		000331 => x"c0a2", -- LDIL
		000332 => x"bee2", -- BL
		000333 => x"24a2", -- LDUB
		000334 => x"3c90", -- SFT
		000335 => x"bedf", -- BL
		000336 => x"3c90", -- SFT
		000337 => x"bedd", -- BL
		000338 => x"24b3", -- LDUB
		000339 => x"3c90", -- SFT
		000340 => x"beda", -- BL
		000341 => x"3c90", -- SFT
		000342 => x"bed8", -- BL
		000343 => x"24c4", -- LDUB
		000344 => x"3c90", -- SFT
		000345 => x"bed5", -- BL
		000346 => x"3c90", -- SFT
		000347 => x"bed3", -- BL
		000348 => x"24d5", -- LDUB
		000349 => x"3c90", -- SFT
		000350 => x"bed0", -- BL
		000351 => x"3c90", -- SFT
		000352 => x"bece", -- BL
		000353 => x"24e6", -- LDUB
		000354 => x"3c90", -- SFT
		000355 => x"becb", -- BL
		000356 => x"3c90", -- SFT
		000357 => x"bec9", -- BL
		000358 => x"c0a2", -- LDIL
		000359 => x"bec7", -- BL
		000360 => x"bec1", -- BL
		000361 => x"c55a", -- LDIL
		000362 => x"c906", -- LDIH
		000363 => x"beb1", -- BL
		000364 => x"2677", -- LDUB
		000365 => x"be4e", -- BL
		000366 => x"bebb", -- BL
		000367 => x"beba", -- BL
		000368 => x"2800", -- CLR
		000369 => x"d58e", -- SBR
		000370 => x"d5bf", -- SBR
		000371 => x"1c03", -- STSR
		000372 => x"ed0f", -- MCR
		000373 => x"ec88", -- MCR
		000374 => x"ec8b", -- MCR
		000375 => x"ec8c", -- MCR
		000376 => x"ec8a", -- MCR
		000377 => x"ec89", -- MCR
		000378 => x"3400", -- GT
		000379 => x"c544", -- LDIL
		000380 => x"c906", -- LDIH
		000381 => x"be9f", -- BL
		000382 => x"beba", -- BL
		000383 => x"beb4", -- BL
		000384 => x"c08d", -- LDIL
		000385 => x"1809", -- CMP
		000386 => x"8006", -- BEQ
		000387 => x"c088", -- LDIL
		000388 => x"1809", -- CMP
		000389 => x"85fa", -- BNE
		000390 => x"bea3", -- BL
		000391 => x"bdbd", -- B
		000392 => x"ecca", -- MCR
		000393 => x"bea0", -- BL
		000394 => x"c280", -- LDIL
		000395 => x"c00f", -- LDIL
		000396 => x"2058", -- ANDS
		000397 => x"840a", -- BNE
		000398 => x"be9b", -- BL
		000399 => x"c0a4", -- LDIL
		000400 => x"be9e", -- BL
		000401 => x"0250", -- MOV
		000402 => x"becb", -- BL
		000403 => x"c0ba", -- LDIL
		000404 => x"be9a", -- BL
		000405 => x"c0a0", -- LDIL
		000406 => x"be98", -- BL
		000407 => x"7a5a", -- LDR
		000408 => x"c0a0", -- LDIL
		000409 => x"be95", -- BL
		000410 => x"bec3", -- BL
		000411 => x"c00f", -- LDIL
		000412 => x"2058", -- ANDS
		000413 => x"8414", -- BNE
		000414 => x"c0a0", -- LDIL
		000415 => x"be8f", -- BL
		000416 => x"be8e", -- BL
		000417 => x"c010", -- LDIL
		000418 => x"1250", -- SUB
		000419 => x"c470", -- LDIL
		000420 => x"2240", -- AND
		000421 => x"78c9", -- LDR
		000422 => x"3c90", -- SFT
		000423 => x"c880", -- LDIH
		000424 => x"c020", -- LDIL
		000425 => x"1818", -- CMP
		000426 => x"a402", -- BLS
		000427 => x"c0ae", -- LDIL
		000428 => x"be82", -- BL
		000429 => x"c08f", -- LDIL
		000430 => x"2014", -- AND
		000431 => x"3409", -- TEQ
		000432 => x"85f5", -- BNE
		000433 => x"ec20", -- MRC
		000434 => x"dc0f", -- STB
		000435 => x"b804", -- BTS
		000436 => x"c5fe", -- LDIL
		000437 => x"343d", -- TEQ
		000438 => x"85d5", -- BNE
		000439 => x"be7c", -- BL
		000440 => x"2800", -- CLR
		000441 => x"3400", -- GT
		000442 => x"bc5e", -- B
		000443 => x"bca2", -- B
		000444 => x"c001", -- LDIL
		000445 => x"ed0c", -- MCR
		000446 => x"c050", -- LDIL
		000447 => x"c83f", -- LDIH
		000448 => x"ed0a", -- MCR
		000449 => x"c000", -- LDIL
		000450 => x"c801", -- LDIH
		000451 => x"beb8", -- BL
		000452 => x"c15e", -- LDIL
		000453 => x"c906", -- LDIH
		000454 => x"be53", -- BL
		000455 => x"c16e", -- LDIL
		000456 => x"c906", -- LDIH
		000457 => x"be50", -- BL
		000458 => x"be69", -- BL
		000459 => x"3c80", -- SFT
		000460 => x"be67", -- BL
		000461 => x"2410", -- ORR
		000462 => x"c4fe", -- LDIL
		000463 => x"ccca", -- LDIH
		000464 => x"1809", -- CMP
		000465 => x"843e", -- BNE
		000466 => x"c100", -- LDIL
		000467 => x"c5ca", -- LDIL
		000468 => x"bead", -- BL
		000469 => x"c101", -- LDIL
		000470 => x"c5fe", -- LDIL
		000471 => x"beaa", -- BL
		000472 => x"be5b", -- BL
		000473 => x"3c80", -- SFT
		000474 => x"be59", -- BL
		000475 => x"2690", -- ORR
		000476 => x"3ed4", -- SFT
		000477 => x"2055", -- STUB
		000478 => x"c102", -- LDIL
		000479 => x"3dd0", -- SFT
		000480 => x"bea1", -- BL
		000481 => x"c103", -- LDIL
		000482 => x"01d0", -- MOV
		000483 => x"be9e", -- BL
		000484 => x"be4f", -- BL
		000485 => x"3c80", -- SFT
		000486 => x"be4d", -- BL
		000487 => x"2690", -- ORR
		000488 => x"20d5", -- STUB
		000489 => x"c104", -- LDIL
		000490 => x"3dd0", -- SFT
		000491 => x"be96", -- BL
		000492 => x"c105", -- LDIL
		000493 => x"01d0", -- MOV
		000494 => x"be93", -- BL
		000495 => x"c106", -- LDIL
		000496 => x"be43", -- BL
		000497 => x"0180", -- MOV
		000498 => x"be8f", -- BL
		000499 => x"0121", -- INC
		000500 => x"c010", -- LDIL
		000501 => x"1828", -- CMP
		000502 => x"85fa", -- BNE
		000503 => x"c110", -- LDIL
		000504 => x"2ad5", -- CLR
		000505 => x"be3a", -- BL
		000506 => x"0180", -- MOV
		000507 => x"be86", -- BL
		000508 => x"0121", -- INC
		000509 => x"2400", -- LDUB
		000510 => x"02d1", -- INC
		000511 => x"1858", -- CMP
		000512 => x"85f9", -- BNE
		000513 => x"c001", -- LDIL
		000514 => x"ed0c", -- MCR
		000515 => x"c050", -- LDIL
		000516 => x"c83f", -- LDIH
		000517 => x"ed0a", -- MCR
		000518 => x"c00c", -- LDIL
		000519 => x"c801", -- LDIH
		000520 => x"be73", -- BL
		000521 => x"c530", -- LDIL
		000522 => x"c906", -- LDIH
		000523 => x"be0e", -- BL
		000524 => x"c6a2", -- LDIL
		000525 => x"ca80", -- LDIH
		000526 => x"3450", -- GT
		000527 => x"c516", -- LDIL
		000528 => x"c907", -- LDIH
		000529 => x"be08", -- BL
		000530 => x"c552", -- LDIL
		000531 => x"c907", -- LDIH
		000532 => x"be05", -- BL
		000533 => x"be1e", -- BL
		000534 => x"2800", -- CLR
		000535 => x"3400", -- GT
		000536 => x"bc9e", -- B
		000537 => x"c5ff", -- LDIL
		000538 => x"0270", -- MOV
		000539 => x"bc03", -- B
		000540 => x"29b3", -- CLR
		000541 => x"0270", -- MOV
		000542 => x"7829", -- LDR
		000543 => x"c080", -- LDIL
		000544 => x"ccff", -- LDIH
		000545 => x"2081", -- AND
		000546 => x"3c98", -- SFTS
		000547 => x"8003", -- BEQ
		000548 => x"be0a", -- BL
		000549 => x"bdf9", -- B
		000550 => x"03c0", -- MOV
		000551 => x"343b", -- TEQ
		000552 => x"f707", -- RBAEQ
		000553 => x"0170", -- MOV
		000554 => x"c08d", -- LDIL
		000555 => x"be03", -- BL
		000556 => x"c08a", -- LDIL
		000557 => x"03a0", -- MOV
		000558 => x"ec22", -- MRC
		000559 => x"dc05", -- STB
		000560 => x"b9fe", -- BTS
		000561 => x"ed18", -- MCR
		000562 => x"3470", -- RET
		000563 => x"ec20", -- MRC
		000564 => x"dc8f", -- STBI
		000565 => x"b9fe", -- BTS
		000566 => x"c800", -- LDIH
		000567 => x"3470", -- RET
		000568 => x"0170", -- MOV
		000569 => x"c200", -- LDIL
		000570 => x"c184", -- LDIL
		000571 => x"bff8", -- BL
		000572 => x"c0c6", -- LDIL
		000573 => x"1809", -- CMP
		000574 => x"9003", -- BMI
		000575 => x"c0a0", -- LDIL
		000576 => x"1001", -- SUB
		000577 => x"c0b0", -- LDIL
		000578 => x"1809", -- CMP
		000579 => x"91f8", -- BMI
		000580 => x"c0c6", -- LDIL
		000581 => x"1818", -- CMP
		000582 => x"91f5", -- BMI
		000583 => x"c0b9", -- LDIL
		000584 => x"1818", -- CMP
		000585 => x"a404", -- BLS
		000586 => x"c0c1", -- LDIL
		000587 => x"1809", -- CMP
		000588 => x"a1ef", -- BHI
		000589 => x"0080", -- MOV
		000590 => x"bfe0", -- BL
		000591 => x"c030", -- LDIL
		000592 => x"1090", -- SUB
		000593 => x"c009", -- LDIL
		000594 => x"1809", -- CMP
		000595 => x"a402", -- BLS
		000596 => x"0497", -- DEC
		000597 => x"3e42", -- SFT
		000598 => x"3e42", -- SFT
		000599 => x"3e42", -- SFT
		000600 => x"3e42", -- SFT
		000601 => x"2641", -- ORR
		000602 => x"05b9", -- DECS
		000603 => x"85e0", -- BNE
		000604 => x"3420", -- RET
		000605 => x"0370", -- MOV
		000606 => x"3d42", -- SFT
		000607 => x"3d22", -- SFT
		000608 => x"3d22", -- SFT
		000609 => x"3d22", -- SFT
		000610 => x"be0f", -- BL
		000611 => x"bfcb", -- BL
		000612 => x"3d40", -- SFT
		000613 => x"be0c", -- BL
		000614 => x"bfc8", -- BL
		000615 => x"3d45", -- SFT
		000616 => x"3d25", -- SFT
		000617 => x"3d25", -- SFT
		000618 => x"3d25", -- SFT
		000619 => x"be06", -- BL
		000620 => x"bfc2", -- BL
		000621 => x"0140", -- MOV
		000622 => x"be03", -- BL
		000623 => x"bfbf", -- BL
		000624 => x"3460", -- RET
		000625 => x"c08f", -- LDIL
		000626 => x"2121", -- AND
		000627 => x"c089", -- LDIL
		000628 => x"181a", -- CMP
		000629 => x"8803", -- BCS
		000630 => x"c0b0", -- LDIL
		000631 => x"bc02", -- B
		000632 => x"c0b7", -- LDIL
		000633 => x"0892", -- ADD
		000634 => x"3470", -- RET
		000635 => x"ed0b", -- MCR
		000636 => x"ec22", -- MRC
		000637 => x"dc03", -- STB
		000638 => x"b9fe", -- BTS
		000639 => x"ec23", -- MRC
		000640 => x"3470", -- RET
		000641 => x"00f0", -- MOV
		000642 => x"c050", -- LDIL
		000643 => x"c837", -- LDIH
		000644 => x"ed0a", -- MCR
		000645 => x"c001", -- LDIL
		000646 => x"ed0c", -- MCR
		000647 => x"c006", -- LDIL
		000648 => x"bff3", -- BL
		000649 => x"c050", -- LDIL
		000650 => x"c83f", -- LDIH
		000651 => x"ed0a", -- MCR
		000652 => x"c000", -- LDIL
		000653 => x"c805", -- LDIH
		000654 => x"bfed", -- BL
		000655 => x"dc01", -- STB
		000656 => x"b80a", -- BTS
		000657 => x"c540", -- LDIL
		000658 => x"c907", -- LDIH
		000659 => x"bf86", -- BL
		000660 => x"c552", -- LDIL
		000661 => x"c907", -- LDIH
		000662 => x"bf83", -- BL
		000663 => x"bf9c", -- BL
		000664 => x"2800", -- CLR
		000665 => x"3400", -- GT
		000666 => x"c040", -- LDIL
		000667 => x"c83f", -- LDIH
		000668 => x"ed0a", -- MCR
		000669 => x"c001", -- LDIL
		000670 => x"ed0c", -- MCR
		000671 => x"3c20", -- SFT
		000672 => x"c802", -- LDIH
		000673 => x"bfda", -- BL
		000674 => x"03a0", -- MOV
		000675 => x"cb80", -- LDIH
		000676 => x"3ff0", -- SFT
		000677 => x"0030", -- MOV
		000678 => x"c800", -- LDIH
		000679 => x"2407", -- ORR
		000680 => x"bfd3", -- BL
		000681 => x"2800", -- CLR
		000682 => x"ed0c", -- MCR
		000683 => x"c050", -- LDIL
		000684 => x"c83f", -- LDIH
		000685 => x"ed0a", -- MCR
		000686 => x"c001", -- LDIL
		000687 => x"ed0c", -- MCR
		000688 => x"c000", -- LDIL
		000689 => x"c805", -- LDIH
		000690 => x"bfc9", -- BL
		000691 => x"dc00", -- STB
		000692 => x"b9fc", -- BTS
		000693 => x"3410", -- RET
		000694 => x"00f0", -- MOV
		000695 => x"c040", -- LDIL
		000696 => x"c83f", -- LDIH
		000697 => x"ed0a", -- MCR
		000698 => x"c001", -- LDIL
		000699 => x"ed0c", -- MCR
		000700 => x"3c20", -- SFT
		000701 => x"c803", -- LDIH
		000702 => x"bfbd", -- BL
		000703 => x"0020", -- MOV
		000704 => x"c800", -- LDIH
		000705 => x"3c00", -- SFT
		000706 => x"bfb9", -- BL
		000707 => x"29b3", -- CLR
		000708 => x"ed3c", -- MCR
		000709 => x"0180", -- MOV
		000710 => x"c980", -- LDIH
		000711 => x"3410", -- RET
		000712 => x"4154", -- .DW
		000713 => x"4c41", -- .DW
		000714 => x"532d", -- .DW
		000715 => x"324b", -- .DW
		000716 => x"2042", -- .DW
		000717 => x"6f6f", -- .DW
		000718 => x"746c", -- .DW
		000719 => x"6f61", -- .DW
		000720 => x"6465", -- .DW
		000721 => x"7220", -- .DW
		000722 => x"2d20", -- .DW
		000723 => x"5665", -- .DW
		000724 => x"7273", -- .DW
		000725 => x"696f", -- .DW
		000726 => x"6e20", -- .DW
		000727 => x"3230", -- .DW
		000728 => x"3134", -- .DW
		000729 => x"2e30", -- .DW
		000730 => x"332e", -- .DW
		000731 => x"3038", -- .DW
		000732 => x"0000", -- .DW
		000733 => x"6279", -- .DW
		000734 => x"2053", -- .DW
		000735 => x"7465", -- .DW
		000736 => x"7068", -- .DW
		000737 => x"616e", -- .DW
		000738 => x"204e", -- .DW
		000739 => x"6f6c", -- .DW
		000740 => x"7469", -- .DW
		000741 => x"6e67", -- .DW
		000742 => x"2c20", -- .DW
		000743 => x"7374", -- .DW
		000744 => x"6e6f", -- .DW
		000745 => x"6c74", -- .DW
		000746 => x"696e", -- .DW
		000747 => x"6740", -- .DW
		000748 => x"676d", -- .DW
		000749 => x"6169", -- .DW
		000750 => x"6c2e", -- .DW
		000751 => x"636f", -- .DW
		000752 => x"6d00", -- .DW
		000753 => x"7777", -- .DW
		000754 => x"772e", -- .DW
		000755 => x"6f70", -- .DW
		000756 => x"656e", -- .DW
		000757 => x"636f", -- .DW
		000758 => x"7265", -- .DW
		000759 => x"732e", -- .DW
		000760 => x"6f72", -- .DW
		000761 => x"672f", -- .DW
		000762 => x"7072", -- .DW
		000763 => x"6f6a", -- .DW
		000764 => x"6563", -- .DW
		000765 => x"742c", -- .DW
		000766 => x"6174", -- .DW
		000767 => x"6c61", -- .DW
		000768 => x"735f", -- .DW
		000769 => x"636f", -- .DW
		000770 => x"7265", -- .DW
		000771 => x"0000", -- .DW
		000772 => x"426f", -- .DW
		000773 => x"6f74", -- .DW
		000774 => x"6c6f", -- .DW
		000775 => x"6164", -- .DW
		000776 => x"6572", -- .DW
		000777 => x"2073", -- .DW
		000778 => x"7461", -- .DW
		000779 => x"7274", -- .DW
		000780 => x"3a20", -- .DW
		000781 => x"3078", -- .DW
		000782 => x"0000", -- .DW
		000783 => x"436c", -- .DW
		000784 => x"6f63", -- .DW
		000785 => x"6b20", -- .DW
		000786 => x"7370", -- .DW
		000787 => x"6565", -- .DW
		000788 => x"6420", -- .DW
		000789 => x"2848", -- .DW
		000790 => x"7a29", -- .DW
		000791 => x"3a20", -- .DW
		000792 => x"3078", -- .DW
		000793 => x"0000", -- .DW
		000794 => x"426f", -- .DW
		000795 => x"6f74", -- .DW
		000796 => x"696e", -- .DW
		000797 => x"6720", -- .DW
		000798 => x"6672", -- .DW
		000799 => x"6f6d", -- .DW
		000800 => x"2053", -- .DW
		000801 => x"5049", -- .DW
		000802 => x"2045", -- .DW
		000803 => x"4550", -- .DW
		000804 => x"524f", -- .DW
		000805 => x"4d00", -- .DW
		000806 => x"426f", -- .DW
		000807 => x"6f74", -- .DW
		000808 => x"696e", -- .DW
		000809 => x"6720", -- .DW
		000810 => x"6672", -- .DW
		000811 => x"6f6d", -- .DW
		000812 => x"2055", -- .DW
		000813 => x"4152", -- .DW
		000814 => x"5400", -- .DW
		000815 => x"4275", -- .DW
		000816 => x"726e", -- .DW
		000817 => x"696e", -- .DW
		000818 => x"6720", -- .DW
		000819 => x"4545", -- .DW
		000820 => x"5052", -- .DW
		000821 => x"4f4d", -- .DW
		000822 => x"0000", -- .DW
		000823 => x"5761", -- .DW
		000824 => x"6974", -- .DW
		000825 => x"696e", -- .DW
		000826 => x"6720", -- .DW
		000827 => x"666f", -- .DW
		000828 => x"7220", -- .DW
		000829 => x"696d", -- .DW
		000830 => x"6167", -- .DW
		000831 => x"6520", -- .DW
		000832 => x"6461", -- .DW
		000833 => x"7461", -- .DW
		000834 => x"2e2e", -- .DW
		000835 => x"2e00", -- .DW
		000836 => x"426f", -- .DW
		000837 => x"6f74", -- .DW
		000838 => x"696e", -- .DW
		000839 => x"6720", -- .DW
		000840 => x"6672", -- .DW
		000841 => x"6f6d", -- .DW
		000842 => x"206d", -- .DW
		000843 => x"656d", -- .DW
		000844 => x"6f72", -- .DW
		000845 => x"792e", -- .DW
		000846 => x"2e2e", -- .DW
		000847 => x"0000", -- .DW
		000848 => x"5374", -- .DW
		000849 => x"6172", -- .DW
		000850 => x"7469", -- .DW
		000851 => x"6e67", -- .DW
		000852 => x"2069", -- .DW
		000853 => x"6d61", -- .DW
		000854 => x"6765", -- .DW
		000855 => x"2000", -- .DW
		000856 => x"446f", -- .DW
		000857 => x"776e", -- .DW
		000858 => x"6c6f", -- .DW
		000859 => x"6164", -- .DW
		000860 => x"2063", -- .DW
		000861 => x"6f6d", -- .DW
		000862 => x"706c", -- .DW
		000863 => x"6574", -- .DW
		000864 => x"6564", -- .DW
		000865 => x"2100", -- .DW
		000866 => x"456e", -- .DW
		000867 => x"7465", -- .DW
		000868 => x"7220", -- .DW
		000869 => x"7061", -- .DW
		000870 => x"6765", -- .DW
		000871 => x"2028", -- .DW
		000872 => x"3468", -- .DW
		000873 => x"6578", -- .DW
		000874 => x"293a", -- .DW
		000875 => x"2030", -- .DW
		000876 => x"7800", -- .DW
		000877 => x"4368", -- .DW
		000878 => x"6563", -- .DW
		000879 => x"6b73", -- .DW
		000880 => x"756d", -- .DW
		000881 => x"3a20", -- .DW
		000882 => x"3078", -- .DW
		000883 => x"0000", -- .DW
		000884 => x"436f", -- .DW
		000885 => x"6d6d", -- .DW
		000886 => x"616e", -- .DW
		000887 => x"642f", -- .DW
		000888 => x"626f", -- .DW
		000889 => x"6f74", -- .DW
		000890 => x"2073", -- .DW
		000891 => x"7769", -- .DW
		000892 => x"7463", -- .DW
		000893 => x"6800", -- .DW
		000894 => x"2030", -- .DW
		000895 => x"2f27", -- .DW
		000896 => x"3030", -- .DW
		000897 => x"273a", -- .DW
		000898 => x"2052", -- .DW
		000899 => x"6573", -- .DW
		000900 => x"7461", -- .DW
		000901 => x"7274", -- .DW
		000902 => x"2063", -- .DW
		000903 => x"6f6e", -- .DW
		000904 => x"736f", -- .DW
		000905 => x"6c65", -- .DW
		000906 => x"0000", -- .DW
		000907 => x"2031", -- .DW
		000908 => x"2f27", -- .DW
		000909 => x"3031", -- .DW
		000910 => x"273a", -- .DW
		000911 => x"2042", -- .DW
		000912 => x"6f6f", -- .DW
		000913 => x"7420", -- .DW
		000914 => x"6672", -- .DW
		000915 => x"6f6d", -- .DW
		000916 => x"2055", -- .DW
		000917 => x"4152", -- .DW
		000918 => x"5400", -- .DW
		000919 => x"2032", -- .DW
		000920 => x"2f27", -- .DW
		000921 => x"3130", -- .DW
		000922 => x"273a", -- .DW
		000923 => x"2042", -- .DW
		000924 => x"6f6f", -- .DW
		000925 => x"7420", -- .DW
		000926 => x"6672", -- .DW
		000927 => x"6f6d", -- .DW
		000928 => x"2045", -- .DW
		000929 => x"4550", -- .DW
		000930 => x"524f", -- .DW
		000931 => x"4d00", -- .DW
		000932 => x"2033", -- .DW
		000933 => x"2f27", -- .DW
		000934 => x"3131", -- .DW
		000935 => x"273a", -- .DW
		000936 => x"2042", -- .DW
		000937 => x"6f6f", -- .DW
		000938 => x"7420", -- .DW
		000939 => x"6672", -- .DW
		000940 => x"6f6d", -- .DW
		000941 => x"206d", -- .DW
		000942 => x"656d", -- .DW
		000943 => x"6f72", -- .DW
		000944 => x"7900", -- .DW
		000945 => x"2070", -- .DW
		000946 => x"3a20", -- .DW
		000947 => x"5072", -- .DW
		000948 => x"6f67", -- .DW
		000949 => x"7261", -- .DW
		000950 => x"6d20", -- .DW
		000951 => x"4545", -- .DW
		000952 => x"5052", -- .DW
		000953 => x"4f4d", -- .DW
		000954 => x"0000", -- .DW
		000955 => x"2064", -- .DW
		000956 => x"3a20", -- .DW
		000957 => x"5241", -- .DW
		000958 => x"4d20", -- .DW
		000959 => x"6475", -- .DW
		000960 => x"6d70", -- .DW
		000961 => x"0000", -- .DW
		000962 => x"2072", -- .DW
		000963 => x"3a20", -- .DW
		000964 => x"5265", -- .DW
		000965 => x"7365", -- .DW
		000966 => x"7400", -- .DW
		000967 => x"636d", -- .DW
		000968 => x"643a", -- .DW
		000969 => x"3e20", -- .DW
		000970 => x"0000", -- .DW
		000971 => x"494d", -- .DW
		000972 => x"4147", -- .DW
		000973 => x"4520", -- .DW
		000974 => x"4552", -- .DW
		000975 => x"524f", -- .DW
		000976 => x"5221", -- .DW
		000977 => x"0000", -- .DW
		000978 => x"4952", -- .DW
		000979 => x"5120", -- .DW
		000980 => x"4552", -- .DW
		000981 => x"524f", -- .DW
		000982 => x"5221", -- .DW
		000983 => x"0000", -- .DW
		000984 => x"4348", -- .DW
		000985 => x"4543", -- .DW
		000986 => x"4b53", -- .DW
		000987 => x"554d", -- .DW
		000988 => x"2045", -- .DW
		000989 => x"5252", -- .DW
		000990 => x"4f52", -- .DW
		000991 => x"2100", -- .DW
		000992 => x"5350", -- .DW
		000993 => x"492f", -- .DW
		000994 => x"4545", -- .DW
		000995 => x"5052", -- .DW
		000996 => x"4f4d", -- .DW
		000997 => x"2045", -- .DW
		000998 => x"5252", -- .DW
		000999 => x"4f52", -- .DW
		001000 => x"2100", -- .DW
		001001 => x"5072", -- .DW
		001002 => x"6573", -- .DW
		001003 => x"7320", -- .DW
		001004 => x"616e", -- .DW
		001005 => x"7920", -- .DW
		001006 => x"6b65", -- .DW
		001007 => x"7900", -- .DW
		others => x"0000"  -- NOP
	);
	------------------------------------------------------

begin

	-- Memory Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		MEM_FILE_ACCESS: process(CLK_I)
		begin
			if rising_edge(CLK_I) then
				-- Data Read --
				if (D_EN_I = '1') then -- valid access
					if (word_mode_en_c = true) then -- read data access
						D_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(D_ADR_I(log2_mem_size_c-1 downto 0))));
					else
						D_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(D_ADR_I(log2_mem_size_c downto 1))));
					end if;
				end if;
				-- Instruction Read --
				if (I_EN_I = '1') then
					if (word_mode_en_c = true) then
						I_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(I_ADR_I(log2_mem_size_c-1 downto 0))));
					else
						I_DAT_O <= BOOT_MEM_FILE_C(to_integer(unsigned(I_ADR_I(log2_mem_size_c downto 1))));
					end if;
				end if;
			end if;
		end process MEM_FILE_ACCESS;



end BOOT_MEM_STRUCTURE;
