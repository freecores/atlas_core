000000 => x"cafe",
000001 => x"00be",
000002 => x"7740",
000003 => x"5241",
000004 => x"4e44",
000005 => x"4f4d",
000006 => x"5f4e",
000007 => x"554d",
000008 => x"bc0b",
000009 => x"bc04",
000010 => x"bc03",
000011 => x"bc02",
000012 => x"bc01",
000013 => x"be31",
000014 => x"c110",
000015 => x"c901",
000016 => x"be21",
000017 => x"be2d",
000018 => x"bc00",
000019 => x"c12c",
000020 => x"c901",
000021 => x"be19",
000022 => x"c144",
000023 => x"c901",
000024 => x"be19",
000025 => x"be34",
000026 => x"ec4d",
000027 => x"be23",
000028 => x"c160",
000029 => x"c901",
000030 => x"be13",
000031 => x"be2e",
000032 => x"d24f",
000033 => x"ec4e",
000034 => x"be1c",
000035 => x"c0b0",
000036 => x"be1f",
000037 => x"c0f8",
000038 => x"be1d",
000039 => x"ee05",
000040 => x"be4a",
000041 => x"be15",
000042 => x"ec20",
000043 => x"dc0f",
000044 => x"b9ea",
000045 => x"bdf6",
000046 => x"c5ff",
000047 => x"0270",
000048 => x"bc03",
000049 => x"29b3",
000050 => x"0270",
000051 => x"7829",
000052 => x"c080",
000053 => x"ccff",
000054 => x"2081",
000055 => x"3c98",
000056 => x"8003",
000057 => x"be0a",
000058 => x"bdf9",
000059 => x"03c0",
000060 => x"343b",
000061 => x"f707",
000062 => x"0170",
000063 => x"c08d",
000064 => x"be03",
000065 => x"c08a",
000066 => x"03a0",
000067 => x"ec22",
000068 => x"dc05",
000069 => x"b9fe",
000070 => x"ed18",
000071 => x"3470",
000072 => x"ec20",
000073 => x"dc8f",
000074 => x"b9fe",
000075 => x"c800",
000076 => x"3470",
000077 => x"0170",
000078 => x"c200",
000079 => x"c184",
000080 => x"bff8",
000081 => x"c0c6",
000082 => x"1809",
000083 => x"9003",
000084 => x"c0a0",
000085 => x"1001",
000086 => x"c0b0",
000087 => x"1809",
000088 => x"91f8",
000089 => x"c0c6",
000090 => x"1818",
000091 => x"91f5",
000092 => x"c0b9",
000093 => x"1818",
000094 => x"a404",
000095 => x"c0c1",
000096 => x"1809",
000097 => x"a1ef",
000098 => x"0080",
000099 => x"bfe0",
000100 => x"c030",
000101 => x"1090",
000102 => x"c009",
000103 => x"1809",
000104 => x"a402",
000105 => x"0497",
000106 => x"3e42",
000107 => x"3e42",
000108 => x"3e42",
000109 => x"3e42",
000110 => x"2641",
000111 => x"05b9",
000112 => x"85e0",
000113 => x"3420",
000114 => x"0370",
000115 => x"3d42",
000116 => x"3d22",
000117 => x"3d22",
000118 => x"3d22",
000119 => x"be0f",
000120 => x"bfcb",
000121 => x"3d40",
000122 => x"be0c",
000123 => x"bfc8",
000124 => x"3d45",
000125 => x"3d25",
000126 => x"3d25",
000127 => x"3d25",
000128 => x"be06",
000129 => x"bfc2",
000130 => x"0140",
000131 => x"be03",
000132 => x"bfbf",
000133 => x"3460",
000134 => x"c08f",
000135 => x"2121",
000136 => x"c089",
000137 => x"181a",
000138 => x"8803",
000139 => x"c0b0",
000140 => x"bc02",
000141 => x"c0b7",
000142 => x"0892",
000143 => x"3470",
000144 => x"4578",
000145 => x"6365",
000146 => x"7074",
000147 => x"696f",
000148 => x"6e2f",
000149 => x"696e",
000150 => x"7465",
000151 => x"7272",
000152 => x"7570",
000153 => x"7420",
000154 => x"6572",
000155 => x"726f",
000156 => x"7221",
000157 => x"0000",
000158 => x"5261",
000159 => x"6e64",
000160 => x"6f6d",
000161 => x"204e",
000162 => x"756d",
000163 => x"6265",
000164 => x"7220",
000165 => x"4765",
000166 => x"6e65",
000167 => x"7261",
000168 => x"746f",
000169 => x"7200",
000170 => x"456e",
000171 => x"7465",
000172 => x"7220",
000173 => x"4c46",
000174 => x"5352",
000175 => x"2073",
000176 => x"6565",
000177 => x"6420",
000178 => x"2834",
000179 => x"6865",
000180 => x"7829",
000181 => x"3a20",
000182 => x"3078",
000183 => x"0000",
000184 => x"456e",
000185 => x"7465",
000186 => x"7220",
000187 => x"4c46",
000188 => x"5352",
000189 => x"2074",
000190 => x"6170",
000191 => x"7320",
000192 => x"2834",
000193 => x"6865",
000194 => x"7829",
000195 => x"3a20",
000196 => x"3078",
000197 => x"0000",
others => x"0000"